// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"
// CREATED		"Fri Mar 24 16:56:27 2023"

module Multiplier_32(
	A,
	B,
	Z
);


input wire	[31:0] A;
input wire	[31:0] B;
output wire	[63:0] Z;

wire	[63:0] Z_ALTERA_SYNTHESIZED;
wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_19;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_25;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_30;
wire	SYNTHESIZED_WIRE_31;
wire	SYNTHESIZED_WIRE_32;
wire	SYNTHESIZED_WIRE_33;
wire	SYNTHESIZED_WIRE_34;
wire	SYNTHESIZED_WIRE_35;
wire	SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_38;
wire	SYNTHESIZED_WIRE_39;
wire	SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_41;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_45;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_47;
wire	SYNTHESIZED_WIRE_48;
wire	SYNTHESIZED_WIRE_49;
wire	SYNTHESIZED_WIRE_50;
wire	SYNTHESIZED_WIRE_51;
wire	SYNTHESIZED_WIRE_52;
wire	SYNTHESIZED_WIRE_53;
wire	SYNTHESIZED_WIRE_54;
wire	SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_57;
wire	SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_60;
wire	SYNTHESIZED_WIRE_61;
wire	SYNTHESIZED_WIRE_62;
wire	SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_66;
wire	SYNTHESIZED_WIRE_67;
wire	SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_69;
wire	SYNTHESIZED_WIRE_70;
wire	SYNTHESIZED_WIRE_71;
wire	SYNTHESIZED_WIRE_72;
wire	SYNTHESIZED_WIRE_73;
wire	SYNTHESIZED_WIRE_74;
wire	SYNTHESIZED_WIRE_75;
wire	SYNTHESIZED_WIRE_76;
wire	SYNTHESIZED_WIRE_77;
wire	SYNTHESIZED_WIRE_78;
wire	SYNTHESIZED_WIRE_79;
wire	SYNTHESIZED_WIRE_80;
wire	SYNTHESIZED_WIRE_81;
wire	SYNTHESIZED_WIRE_82;
wire	SYNTHESIZED_WIRE_83;
wire	SYNTHESIZED_WIRE_84;
wire	SYNTHESIZED_WIRE_85;
wire	SYNTHESIZED_WIRE_86;
wire	SYNTHESIZED_WIRE_87;
wire	SYNTHESIZED_WIRE_88;
wire	SYNTHESIZED_WIRE_89;
wire	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_91;
wire	SYNTHESIZED_WIRE_92;
wire	SYNTHESIZED_WIRE_93;
wire	SYNTHESIZED_WIRE_94;
wire	SYNTHESIZED_WIRE_95;
wire	SYNTHESIZED_WIRE_96;
wire	SYNTHESIZED_WIRE_97;
wire	SYNTHESIZED_WIRE_98;
wire	SYNTHESIZED_WIRE_99;
wire	SYNTHESIZED_WIRE_100;
wire	SYNTHESIZED_WIRE_101;
wire	SYNTHESIZED_WIRE_102;
wire	SYNTHESIZED_WIRE_103;
wire	SYNTHESIZED_WIRE_104;
wire	SYNTHESIZED_WIRE_105;
wire	SYNTHESIZED_WIRE_106;
wire	SYNTHESIZED_WIRE_107;
wire	SYNTHESIZED_WIRE_108;
wire	SYNTHESIZED_WIRE_109;
wire	SYNTHESIZED_WIRE_110;
wire	SYNTHESIZED_WIRE_111;
wire	SYNTHESIZED_WIRE_112;
wire	SYNTHESIZED_WIRE_113;
wire	SYNTHESIZED_WIRE_114;
wire	SYNTHESIZED_WIRE_115;
wire	SYNTHESIZED_WIRE_116;
wire	SYNTHESIZED_WIRE_117;
wire	SYNTHESIZED_WIRE_118;
wire	SYNTHESIZED_WIRE_119;
wire	SYNTHESIZED_WIRE_120;
wire	SYNTHESIZED_WIRE_121;
wire	SYNTHESIZED_WIRE_122;
wire	SYNTHESIZED_WIRE_123;
wire	SYNTHESIZED_WIRE_124;
wire	SYNTHESIZED_WIRE_125;
wire	SYNTHESIZED_WIRE_126;
wire	SYNTHESIZED_WIRE_127;
wire	SYNTHESIZED_WIRE_128;
wire	SYNTHESIZED_WIRE_129;
wire	SYNTHESIZED_WIRE_130;
wire	SYNTHESIZED_WIRE_131;
wire	SYNTHESIZED_WIRE_132;
wire	SYNTHESIZED_WIRE_133;
wire	SYNTHESIZED_WIRE_134;
wire	SYNTHESIZED_WIRE_135;
wire	SYNTHESIZED_WIRE_136;
wire	SYNTHESIZED_WIRE_137;
wire	SYNTHESIZED_WIRE_138;
wire	SYNTHESIZED_WIRE_139;
wire	SYNTHESIZED_WIRE_140;
wire	SYNTHESIZED_WIRE_141;
wire	SYNTHESIZED_WIRE_142;
wire	SYNTHESIZED_WIRE_143;
wire	SYNTHESIZED_WIRE_144;
wire	SYNTHESIZED_WIRE_145;
wire	SYNTHESIZED_WIRE_146;
wire	SYNTHESIZED_WIRE_147;
wire	SYNTHESIZED_WIRE_148;
wire	SYNTHESIZED_WIRE_149;
wire	SYNTHESIZED_WIRE_150;
wire	SYNTHESIZED_WIRE_151;
wire	SYNTHESIZED_WIRE_152;
wire	SYNTHESIZED_WIRE_153;
wire	SYNTHESIZED_WIRE_154;
wire	SYNTHESIZED_WIRE_155;
wire	SYNTHESIZED_WIRE_156;
wire	SYNTHESIZED_WIRE_157;
wire	SYNTHESIZED_WIRE_158;
wire	SYNTHESIZED_WIRE_159;
wire	SYNTHESIZED_WIRE_160;
wire	SYNTHESIZED_WIRE_161;
wire	SYNTHESIZED_WIRE_162;
wire	SYNTHESIZED_WIRE_163;
wire	SYNTHESIZED_WIRE_164;
wire	SYNTHESIZED_WIRE_165;
wire	SYNTHESIZED_WIRE_166;
wire	SYNTHESIZED_WIRE_167;
wire	SYNTHESIZED_WIRE_168;
wire	SYNTHESIZED_WIRE_169;
wire	SYNTHESIZED_WIRE_170;
wire	SYNTHESIZED_WIRE_171;
wire	SYNTHESIZED_WIRE_172;
wire	SYNTHESIZED_WIRE_173;
wire	SYNTHESIZED_WIRE_174;
wire	SYNTHESIZED_WIRE_175;
wire	SYNTHESIZED_WIRE_176;
wire	SYNTHESIZED_WIRE_177;
wire	SYNTHESIZED_WIRE_178;
wire	SYNTHESIZED_WIRE_179;
wire	SYNTHESIZED_WIRE_180;
wire	SYNTHESIZED_WIRE_181;
wire	SYNTHESIZED_WIRE_182;
wire	SYNTHESIZED_WIRE_183;
wire	SYNTHESIZED_WIRE_184;
wire	SYNTHESIZED_WIRE_185;
wire	SYNTHESIZED_WIRE_186;
wire	SYNTHESIZED_WIRE_187;
wire	SYNTHESIZED_WIRE_188;
wire	SYNTHESIZED_WIRE_189;
wire	SYNTHESIZED_WIRE_190;
wire	SYNTHESIZED_WIRE_191;
wire	SYNTHESIZED_WIRE_192;
wire	SYNTHESIZED_WIRE_193;
wire	SYNTHESIZED_WIRE_194;
wire	SYNTHESIZED_WIRE_195;
wire	SYNTHESIZED_WIRE_196;
wire	SYNTHESIZED_WIRE_197;
wire	SYNTHESIZED_WIRE_198;
wire	SYNTHESIZED_WIRE_199;
wire	SYNTHESIZED_WIRE_200;
wire	SYNTHESIZED_WIRE_201;
wire	SYNTHESIZED_WIRE_202;
wire	SYNTHESIZED_WIRE_203;
wire	SYNTHESIZED_WIRE_204;
wire	SYNTHESIZED_WIRE_205;
wire	SYNTHESIZED_WIRE_206;
wire	SYNTHESIZED_WIRE_207;
wire	SYNTHESIZED_WIRE_208;
wire	SYNTHESIZED_WIRE_209;
wire	SYNTHESIZED_WIRE_210;
wire	SYNTHESIZED_WIRE_211;
wire	SYNTHESIZED_WIRE_212;
wire	SYNTHESIZED_WIRE_213;
wire	SYNTHESIZED_WIRE_214;
wire	SYNTHESIZED_WIRE_215;
wire	SYNTHESIZED_WIRE_216;
wire	SYNTHESIZED_WIRE_217;
wire	SYNTHESIZED_WIRE_218;
wire	SYNTHESIZED_WIRE_219;
wire	SYNTHESIZED_WIRE_220;
wire	SYNTHESIZED_WIRE_221;
wire	SYNTHESIZED_WIRE_222;
wire	SYNTHESIZED_WIRE_223;
wire	SYNTHESIZED_WIRE_224;
wire	SYNTHESIZED_WIRE_225;
wire	SYNTHESIZED_WIRE_226;
wire	SYNTHESIZED_WIRE_227;
wire	SYNTHESIZED_WIRE_228;
wire	SYNTHESIZED_WIRE_229;
wire	SYNTHESIZED_WIRE_230;
wire	SYNTHESIZED_WIRE_231;
wire	SYNTHESIZED_WIRE_232;
wire	SYNTHESIZED_WIRE_233;
wire	SYNTHESIZED_WIRE_234;
wire	SYNTHESIZED_WIRE_235;
wire	SYNTHESIZED_WIRE_236;
wire	SYNTHESIZED_WIRE_237;
wire	SYNTHESIZED_WIRE_238;
wire	SYNTHESIZED_WIRE_239;
wire	SYNTHESIZED_WIRE_240;
wire	SYNTHESIZED_WIRE_241;
wire	SYNTHESIZED_WIRE_242;
wire	SYNTHESIZED_WIRE_243;
wire	SYNTHESIZED_WIRE_244;
wire	SYNTHESIZED_WIRE_245;
wire	SYNTHESIZED_WIRE_246;
wire	SYNTHESIZED_WIRE_247;
wire	SYNTHESIZED_WIRE_248;
wire	SYNTHESIZED_WIRE_249;
wire	SYNTHESIZED_WIRE_250;
wire	SYNTHESIZED_WIRE_251;
wire	SYNTHESIZED_WIRE_252;
wire	SYNTHESIZED_WIRE_253;
wire	SYNTHESIZED_WIRE_254;
wire	SYNTHESIZED_WIRE_255;
wire	SYNTHESIZED_WIRE_256;
wire	SYNTHESIZED_WIRE_257;
wire	SYNTHESIZED_WIRE_258;
wire	SYNTHESIZED_WIRE_259;
wire	SYNTHESIZED_WIRE_260;
wire	SYNTHESIZED_WIRE_261;
wire	SYNTHESIZED_WIRE_262;
wire	SYNTHESIZED_WIRE_263;
wire	SYNTHESIZED_WIRE_264;
wire	SYNTHESIZED_WIRE_265;
wire	SYNTHESIZED_WIRE_266;
wire	SYNTHESIZED_WIRE_267;
wire	SYNTHESIZED_WIRE_268;
wire	SYNTHESIZED_WIRE_269;
wire	SYNTHESIZED_WIRE_270;
wire	SYNTHESIZED_WIRE_271;
wire	SYNTHESIZED_WIRE_272;
wire	SYNTHESIZED_WIRE_273;
wire	SYNTHESIZED_WIRE_274;
wire	SYNTHESIZED_WIRE_275;
wire	SYNTHESIZED_WIRE_276;
wire	SYNTHESIZED_WIRE_277;
wire	SYNTHESIZED_WIRE_278;
wire	SYNTHESIZED_WIRE_279;
wire	SYNTHESIZED_WIRE_280;
wire	SYNTHESIZED_WIRE_281;
wire	SYNTHESIZED_WIRE_282;
wire	SYNTHESIZED_WIRE_283;
wire	SYNTHESIZED_WIRE_284;
wire	SYNTHESIZED_WIRE_285;
wire	SYNTHESIZED_WIRE_286;
wire	SYNTHESIZED_WIRE_287;
wire	SYNTHESIZED_WIRE_288;
wire	SYNTHESIZED_WIRE_289;
wire	SYNTHESIZED_WIRE_290;
wire	SYNTHESIZED_WIRE_291;
wire	SYNTHESIZED_WIRE_292;
wire	SYNTHESIZED_WIRE_293;
wire	SYNTHESIZED_WIRE_294;
wire	SYNTHESIZED_WIRE_295;
wire	SYNTHESIZED_WIRE_296;
wire	SYNTHESIZED_WIRE_297;
wire	SYNTHESIZED_WIRE_298;
wire	SYNTHESIZED_WIRE_299;
wire	SYNTHESIZED_WIRE_300;
wire	SYNTHESIZED_WIRE_301;
wire	SYNTHESIZED_WIRE_302;
wire	SYNTHESIZED_WIRE_303;
wire	SYNTHESIZED_WIRE_304;
wire	SYNTHESIZED_WIRE_305;
wire	SYNTHESIZED_WIRE_306;
wire	SYNTHESIZED_WIRE_307;
wire	SYNTHESIZED_WIRE_308;
wire	SYNTHESIZED_WIRE_309;
wire	SYNTHESIZED_WIRE_310;
wire	SYNTHESIZED_WIRE_311;
wire	SYNTHESIZED_WIRE_312;
wire	SYNTHESIZED_WIRE_313;
wire	SYNTHESIZED_WIRE_314;
wire	SYNTHESIZED_WIRE_315;
wire	SYNTHESIZED_WIRE_316;
wire	SYNTHESIZED_WIRE_317;
wire	SYNTHESIZED_WIRE_318;
wire	SYNTHESIZED_WIRE_319;
wire	SYNTHESIZED_WIRE_320;
wire	SYNTHESIZED_WIRE_321;
wire	SYNTHESIZED_WIRE_322;
wire	SYNTHESIZED_WIRE_323;
wire	SYNTHESIZED_WIRE_324;
wire	SYNTHESIZED_WIRE_325;
wire	SYNTHESIZED_WIRE_326;
wire	SYNTHESIZED_WIRE_327;
wire	SYNTHESIZED_WIRE_328;
wire	SYNTHESIZED_WIRE_329;
wire	SYNTHESIZED_WIRE_330;
wire	SYNTHESIZED_WIRE_331;
wire	SYNTHESIZED_WIRE_332;
wire	SYNTHESIZED_WIRE_333;
wire	SYNTHESIZED_WIRE_334;
wire	SYNTHESIZED_WIRE_335;
wire	SYNTHESIZED_WIRE_336;
wire	SYNTHESIZED_WIRE_337;
wire	SYNTHESIZED_WIRE_338;
wire	SYNTHESIZED_WIRE_339;
wire	SYNTHESIZED_WIRE_340;
wire	SYNTHESIZED_WIRE_341;
wire	SYNTHESIZED_WIRE_342;
wire	SYNTHESIZED_WIRE_343;
wire	SYNTHESIZED_WIRE_344;
wire	SYNTHESIZED_WIRE_345;
wire	SYNTHESIZED_WIRE_346;
wire	SYNTHESIZED_WIRE_347;
wire	SYNTHESIZED_WIRE_348;
wire	SYNTHESIZED_WIRE_349;
wire	SYNTHESIZED_WIRE_350;
wire	SYNTHESIZED_WIRE_351;
wire	SYNTHESIZED_WIRE_352;
wire	SYNTHESIZED_WIRE_353;
wire	SYNTHESIZED_WIRE_354;
wire	SYNTHESIZED_WIRE_355;
wire	SYNTHESIZED_WIRE_356;
wire	SYNTHESIZED_WIRE_357;
wire	SYNTHESIZED_WIRE_358;
wire	SYNTHESIZED_WIRE_359;
wire	SYNTHESIZED_WIRE_360;
wire	SYNTHESIZED_WIRE_361;
wire	SYNTHESIZED_WIRE_362;
wire	SYNTHESIZED_WIRE_363;
wire	SYNTHESIZED_WIRE_364;
wire	SYNTHESIZED_WIRE_365;
wire	SYNTHESIZED_WIRE_366;
wire	SYNTHESIZED_WIRE_367;
wire	SYNTHESIZED_WIRE_368;
wire	SYNTHESIZED_WIRE_369;
wire	SYNTHESIZED_WIRE_370;
wire	SYNTHESIZED_WIRE_371;
wire	SYNTHESIZED_WIRE_372;
wire	SYNTHESIZED_WIRE_373;
wire	SYNTHESIZED_WIRE_374;
wire	SYNTHESIZED_WIRE_375;
wire	SYNTHESIZED_WIRE_376;
wire	SYNTHESIZED_WIRE_377;
wire	SYNTHESIZED_WIRE_378;
wire	SYNTHESIZED_WIRE_379;
wire	SYNTHESIZED_WIRE_380;
wire	SYNTHESIZED_WIRE_381;
wire	SYNTHESIZED_WIRE_382;
wire	SYNTHESIZED_WIRE_383;
wire	SYNTHESIZED_WIRE_384;
wire	SYNTHESIZED_WIRE_385;
wire	SYNTHESIZED_WIRE_386;
wire	SYNTHESIZED_WIRE_387;
wire	SYNTHESIZED_WIRE_388;
wire	SYNTHESIZED_WIRE_389;
wire	SYNTHESIZED_WIRE_390;
wire	SYNTHESIZED_WIRE_391;
wire	SYNTHESIZED_WIRE_392;
wire	SYNTHESIZED_WIRE_393;
wire	SYNTHESIZED_WIRE_394;
wire	SYNTHESIZED_WIRE_395;
wire	SYNTHESIZED_WIRE_396;
wire	SYNTHESIZED_WIRE_397;
wire	SYNTHESIZED_WIRE_398;
wire	SYNTHESIZED_WIRE_399;
wire	SYNTHESIZED_WIRE_400;
wire	SYNTHESIZED_WIRE_401;
wire	SYNTHESIZED_WIRE_402;
wire	SYNTHESIZED_WIRE_403;
wire	SYNTHESIZED_WIRE_404;
wire	SYNTHESIZED_WIRE_405;
wire	SYNTHESIZED_WIRE_406;
wire	SYNTHESIZED_WIRE_407;
wire	SYNTHESIZED_WIRE_408;
wire	SYNTHESIZED_WIRE_409;
wire	SYNTHESIZED_WIRE_410;
wire	SYNTHESIZED_WIRE_411;
wire	SYNTHESIZED_WIRE_412;
wire	SYNTHESIZED_WIRE_413;
wire	SYNTHESIZED_WIRE_414;
wire	SYNTHESIZED_WIRE_415;
wire	SYNTHESIZED_WIRE_416;
wire	SYNTHESIZED_WIRE_417;
wire	SYNTHESIZED_WIRE_418;
wire	SYNTHESIZED_WIRE_419;
wire	SYNTHESIZED_WIRE_420;
wire	SYNTHESIZED_WIRE_421;
wire	SYNTHESIZED_WIRE_422;
wire	SYNTHESIZED_WIRE_423;
wire	SYNTHESIZED_WIRE_424;
wire	SYNTHESIZED_WIRE_425;
wire	SYNTHESIZED_WIRE_426;
wire	SYNTHESIZED_WIRE_427;
wire	SYNTHESIZED_WIRE_428;
wire	SYNTHESIZED_WIRE_429;
wire	SYNTHESIZED_WIRE_430;
wire	SYNTHESIZED_WIRE_431;
wire	SYNTHESIZED_WIRE_432;
wire	SYNTHESIZED_WIRE_433;
wire	SYNTHESIZED_WIRE_434;
wire	SYNTHESIZED_WIRE_435;
wire	SYNTHESIZED_WIRE_436;
wire	SYNTHESIZED_WIRE_437;
wire	SYNTHESIZED_WIRE_438;
wire	SYNTHESIZED_WIRE_439;
wire	SYNTHESIZED_WIRE_440;
wire	SYNTHESIZED_WIRE_441;
wire	SYNTHESIZED_WIRE_442;
wire	SYNTHESIZED_WIRE_443;
wire	SYNTHESIZED_WIRE_444;
wire	SYNTHESIZED_WIRE_445;
wire	SYNTHESIZED_WIRE_446;
wire	SYNTHESIZED_WIRE_447;
wire	SYNTHESIZED_WIRE_448;
wire	SYNTHESIZED_WIRE_449;
wire	SYNTHESIZED_WIRE_450;
wire	SYNTHESIZED_WIRE_451;
wire	SYNTHESIZED_WIRE_452;
wire	SYNTHESIZED_WIRE_453;
wire	SYNTHESIZED_WIRE_454;
wire	SYNTHESIZED_WIRE_455;
wire	SYNTHESIZED_WIRE_456;
wire	SYNTHESIZED_WIRE_457;
wire	SYNTHESIZED_WIRE_458;
wire	SYNTHESIZED_WIRE_459;
wire	SYNTHESIZED_WIRE_460;
wire	SYNTHESIZED_WIRE_461;
wire	SYNTHESIZED_WIRE_462;
wire	SYNTHESIZED_WIRE_463;
wire	SYNTHESIZED_WIRE_464;
wire	SYNTHESIZED_WIRE_465;
wire	SYNTHESIZED_WIRE_466;
wire	SYNTHESIZED_WIRE_467;
wire	SYNTHESIZED_WIRE_468;
wire	SYNTHESIZED_WIRE_469;
wire	SYNTHESIZED_WIRE_470;
wire	SYNTHESIZED_WIRE_471;
wire	SYNTHESIZED_WIRE_472;
wire	SYNTHESIZED_WIRE_473;
wire	SYNTHESIZED_WIRE_474;
wire	SYNTHESIZED_WIRE_475;
wire	SYNTHESIZED_WIRE_476;
wire	SYNTHESIZED_WIRE_477;
wire	SYNTHESIZED_WIRE_478;
wire	SYNTHESIZED_WIRE_479;
wire	SYNTHESIZED_WIRE_480;
wire	SYNTHESIZED_WIRE_481;
wire	SYNTHESIZED_WIRE_482;
wire	SYNTHESIZED_WIRE_483;
wire	SYNTHESIZED_WIRE_484;
wire	SYNTHESIZED_WIRE_485;
wire	SYNTHESIZED_WIRE_486;
wire	SYNTHESIZED_WIRE_487;
wire	SYNTHESIZED_WIRE_488;
wire	SYNTHESIZED_WIRE_489;
wire	SYNTHESIZED_WIRE_490;
wire	SYNTHESIZED_WIRE_491;
wire	SYNTHESIZED_WIRE_492;
wire	SYNTHESIZED_WIRE_493;
wire	SYNTHESIZED_WIRE_494;
wire	SYNTHESIZED_WIRE_495;
wire	SYNTHESIZED_WIRE_496;
wire	SYNTHESIZED_WIRE_497;
wire	SYNTHESIZED_WIRE_498;
wire	SYNTHESIZED_WIRE_499;
wire	SYNTHESIZED_WIRE_500;
wire	SYNTHESIZED_WIRE_501;
wire	SYNTHESIZED_WIRE_502;
wire	SYNTHESIZED_WIRE_503;
wire	SYNTHESIZED_WIRE_504;
wire	SYNTHESIZED_WIRE_505;
wire	SYNTHESIZED_WIRE_506;
wire	SYNTHESIZED_WIRE_507;
wire	SYNTHESIZED_WIRE_508;
wire	SYNTHESIZED_WIRE_509;
wire	SYNTHESIZED_WIRE_510;
wire	SYNTHESIZED_WIRE_511;
wire	SYNTHESIZED_WIRE_512;
wire	SYNTHESIZED_WIRE_513;
wire	SYNTHESIZED_WIRE_514;
wire	SYNTHESIZED_WIRE_515;
wire	SYNTHESIZED_WIRE_516;
wire	SYNTHESIZED_WIRE_517;
wire	SYNTHESIZED_WIRE_518;
wire	SYNTHESIZED_WIRE_519;
wire	SYNTHESIZED_WIRE_520;
wire	SYNTHESIZED_WIRE_521;
wire	SYNTHESIZED_WIRE_522;
wire	SYNTHESIZED_WIRE_523;
wire	SYNTHESIZED_WIRE_524;
wire	SYNTHESIZED_WIRE_525;
wire	SYNTHESIZED_WIRE_526;
wire	SYNTHESIZED_WIRE_527;
wire	SYNTHESIZED_WIRE_528;
wire	SYNTHESIZED_WIRE_529;
wire	SYNTHESIZED_WIRE_530;
wire	SYNTHESIZED_WIRE_531;
wire	SYNTHESIZED_WIRE_532;
wire	SYNTHESIZED_WIRE_533;
wire	SYNTHESIZED_WIRE_534;
wire	SYNTHESIZED_WIRE_535;
wire	SYNTHESIZED_WIRE_536;
wire	SYNTHESIZED_WIRE_537;
wire	SYNTHESIZED_WIRE_538;
wire	SYNTHESIZED_WIRE_539;
wire	SYNTHESIZED_WIRE_540;
wire	SYNTHESIZED_WIRE_541;
wire	SYNTHESIZED_WIRE_542;
wire	SYNTHESIZED_WIRE_543;
wire	SYNTHESIZED_WIRE_544;
wire	SYNTHESIZED_WIRE_545;
wire	SYNTHESIZED_WIRE_546;
wire	SYNTHESIZED_WIRE_547;
wire	SYNTHESIZED_WIRE_548;
wire	SYNTHESIZED_WIRE_549;
wire	SYNTHESIZED_WIRE_550;
wire	SYNTHESIZED_WIRE_551;
wire	SYNTHESIZED_WIRE_552;
wire	SYNTHESIZED_WIRE_553;
wire	SYNTHESIZED_WIRE_554;
wire	SYNTHESIZED_WIRE_555;
wire	SYNTHESIZED_WIRE_556;
wire	SYNTHESIZED_WIRE_557;
wire	SYNTHESIZED_WIRE_558;
wire	SYNTHESIZED_WIRE_559;
wire	SYNTHESIZED_WIRE_560;
wire	SYNTHESIZED_WIRE_561;
wire	SYNTHESIZED_WIRE_562;
wire	SYNTHESIZED_WIRE_563;
wire	SYNTHESIZED_WIRE_564;
wire	SYNTHESIZED_WIRE_565;
wire	SYNTHESIZED_WIRE_566;
wire	SYNTHESIZED_WIRE_567;
wire	SYNTHESIZED_WIRE_568;
wire	SYNTHESIZED_WIRE_569;
wire	SYNTHESIZED_WIRE_570;
wire	SYNTHESIZED_WIRE_571;
wire	SYNTHESIZED_WIRE_572;
wire	SYNTHESIZED_WIRE_573;
wire	SYNTHESIZED_WIRE_574;
wire	SYNTHESIZED_WIRE_575;
wire	SYNTHESIZED_WIRE_576;
wire	SYNTHESIZED_WIRE_577;
wire	SYNTHESIZED_WIRE_578;
wire	SYNTHESIZED_WIRE_579;
wire	SYNTHESIZED_WIRE_580;
wire	SYNTHESIZED_WIRE_581;
wire	SYNTHESIZED_WIRE_582;
wire	SYNTHESIZED_WIRE_583;
wire	SYNTHESIZED_WIRE_584;
wire	SYNTHESIZED_WIRE_585;
wire	SYNTHESIZED_WIRE_586;
wire	SYNTHESIZED_WIRE_587;
wire	SYNTHESIZED_WIRE_588;
wire	SYNTHESIZED_WIRE_589;
wire	SYNTHESIZED_WIRE_590;
wire	SYNTHESIZED_WIRE_591;
wire	SYNTHESIZED_WIRE_592;
wire	SYNTHESIZED_WIRE_593;
wire	SYNTHESIZED_WIRE_594;
wire	SYNTHESIZED_WIRE_595;
wire	SYNTHESIZED_WIRE_596;
wire	SYNTHESIZED_WIRE_597;
wire	SYNTHESIZED_WIRE_598;
wire	SYNTHESIZED_WIRE_599;
wire	SYNTHESIZED_WIRE_600;
wire	SYNTHESIZED_WIRE_601;
wire	SYNTHESIZED_WIRE_602;
wire	SYNTHESIZED_WIRE_603;
wire	SYNTHESIZED_WIRE_604;
wire	SYNTHESIZED_WIRE_605;
wire	SYNTHESIZED_WIRE_606;
wire	SYNTHESIZED_WIRE_607;
wire	SYNTHESIZED_WIRE_608;
wire	SYNTHESIZED_WIRE_609;
wire	SYNTHESIZED_WIRE_610;
wire	SYNTHESIZED_WIRE_611;
wire	SYNTHESIZED_WIRE_612;
wire	SYNTHESIZED_WIRE_613;
wire	SYNTHESIZED_WIRE_614;
wire	SYNTHESIZED_WIRE_615;
wire	SYNTHESIZED_WIRE_616;
wire	SYNTHESIZED_WIRE_617;
wire	SYNTHESIZED_WIRE_618;
wire	SYNTHESIZED_WIRE_619;
wire	SYNTHESIZED_WIRE_620;
wire	SYNTHESIZED_WIRE_621;
wire	SYNTHESIZED_WIRE_622;
wire	SYNTHESIZED_WIRE_623;
wire	SYNTHESIZED_WIRE_624;
wire	SYNTHESIZED_WIRE_625;
wire	SYNTHESIZED_WIRE_626;
wire	SYNTHESIZED_WIRE_627;
wire	SYNTHESIZED_WIRE_628;
wire	SYNTHESIZED_WIRE_629;
wire	SYNTHESIZED_WIRE_630;
wire	SYNTHESIZED_WIRE_631;
wire	SYNTHESIZED_WIRE_632;
wire	SYNTHESIZED_WIRE_633;
wire	SYNTHESIZED_WIRE_634;
wire	SYNTHESIZED_WIRE_635;
wire	SYNTHESIZED_WIRE_636;
wire	SYNTHESIZED_WIRE_637;
wire	SYNTHESIZED_WIRE_638;
wire	SYNTHESIZED_WIRE_639;
wire	SYNTHESIZED_WIRE_640;
wire	SYNTHESIZED_WIRE_641;
wire	SYNTHESIZED_WIRE_642;
wire	SYNTHESIZED_WIRE_643;
wire	SYNTHESIZED_WIRE_644;
wire	SYNTHESIZED_WIRE_645;
wire	SYNTHESIZED_WIRE_646;
wire	SYNTHESIZED_WIRE_647;
wire	SYNTHESIZED_WIRE_648;
wire	SYNTHESIZED_WIRE_649;
wire	SYNTHESIZED_WIRE_650;
wire	SYNTHESIZED_WIRE_651;
wire	SYNTHESIZED_WIRE_652;
wire	SYNTHESIZED_WIRE_653;
wire	SYNTHESIZED_WIRE_654;
wire	SYNTHESIZED_WIRE_655;
wire	SYNTHESIZED_WIRE_656;
wire	SYNTHESIZED_WIRE_657;
wire	SYNTHESIZED_WIRE_658;
wire	SYNTHESIZED_WIRE_659;
wire	SYNTHESIZED_WIRE_660;
wire	SYNTHESIZED_WIRE_661;
wire	SYNTHESIZED_WIRE_662;
wire	SYNTHESIZED_WIRE_663;
wire	SYNTHESIZED_WIRE_664;
wire	SYNTHESIZED_WIRE_665;
wire	SYNTHESIZED_WIRE_666;
wire	SYNTHESIZED_WIRE_667;
wire	SYNTHESIZED_WIRE_668;
wire	SYNTHESIZED_WIRE_669;
wire	SYNTHESIZED_WIRE_670;
wire	SYNTHESIZED_WIRE_671;
wire	SYNTHESIZED_WIRE_672;
wire	SYNTHESIZED_WIRE_673;
wire	SYNTHESIZED_WIRE_674;
wire	SYNTHESIZED_WIRE_675;
wire	SYNTHESIZED_WIRE_676;
wire	SYNTHESIZED_WIRE_677;
wire	SYNTHESIZED_WIRE_678;
wire	SYNTHESIZED_WIRE_679;
wire	SYNTHESIZED_WIRE_680;
wire	SYNTHESIZED_WIRE_681;
wire	SYNTHESIZED_WIRE_682;
wire	SYNTHESIZED_WIRE_683;
wire	SYNTHESIZED_WIRE_684;
wire	SYNTHESIZED_WIRE_685;
wire	SYNTHESIZED_WIRE_686;
wire	SYNTHESIZED_WIRE_687;
wire	SYNTHESIZED_WIRE_688;
wire	SYNTHESIZED_WIRE_689;
wire	SYNTHESIZED_WIRE_690;
wire	SYNTHESIZED_WIRE_691;
wire	SYNTHESIZED_WIRE_692;
wire	SYNTHESIZED_WIRE_693;
wire	SYNTHESIZED_WIRE_694;
wire	SYNTHESIZED_WIRE_695;
wire	SYNTHESIZED_WIRE_696;
wire	SYNTHESIZED_WIRE_697;
wire	SYNTHESIZED_WIRE_698;
wire	SYNTHESIZED_WIRE_699;
wire	SYNTHESIZED_WIRE_700;
wire	SYNTHESIZED_WIRE_701;
wire	SYNTHESIZED_WIRE_702;
wire	SYNTHESIZED_WIRE_703;
wire	SYNTHESIZED_WIRE_704;
wire	SYNTHESIZED_WIRE_705;
wire	SYNTHESIZED_WIRE_706;
wire	SYNTHESIZED_WIRE_707;
wire	SYNTHESIZED_WIRE_708;
wire	SYNTHESIZED_WIRE_709;
wire	SYNTHESIZED_WIRE_710;
wire	SYNTHESIZED_WIRE_711;
wire	SYNTHESIZED_WIRE_712;
wire	SYNTHESIZED_WIRE_713;
wire	SYNTHESIZED_WIRE_714;
wire	SYNTHESIZED_WIRE_715;
wire	SYNTHESIZED_WIRE_716;
wire	SYNTHESIZED_WIRE_717;
wire	SYNTHESIZED_WIRE_718;
wire	SYNTHESIZED_WIRE_719;
wire	SYNTHESIZED_WIRE_720;
wire	SYNTHESIZED_WIRE_721;
wire	SYNTHESIZED_WIRE_722;
wire	SYNTHESIZED_WIRE_723;
wire	SYNTHESIZED_WIRE_724;
wire	SYNTHESIZED_WIRE_725;
wire	SYNTHESIZED_WIRE_726;
wire	SYNTHESIZED_WIRE_727;
wire	SYNTHESIZED_WIRE_728;
wire	SYNTHESIZED_WIRE_729;
wire	SYNTHESIZED_WIRE_730;
wire	SYNTHESIZED_WIRE_731;
wire	SYNTHESIZED_WIRE_732;
wire	SYNTHESIZED_WIRE_733;
wire	SYNTHESIZED_WIRE_734;
wire	SYNTHESIZED_WIRE_735;
wire	SYNTHESIZED_WIRE_736;
wire	SYNTHESIZED_WIRE_737;
wire	SYNTHESIZED_WIRE_738;
wire	SYNTHESIZED_WIRE_739;
wire	SYNTHESIZED_WIRE_740;
wire	SYNTHESIZED_WIRE_741;
wire	SYNTHESIZED_WIRE_742;
wire	SYNTHESIZED_WIRE_743;
wire	SYNTHESIZED_WIRE_744;
wire	SYNTHESIZED_WIRE_745;
wire	SYNTHESIZED_WIRE_746;
wire	SYNTHESIZED_WIRE_747;
wire	SYNTHESIZED_WIRE_748;
wire	SYNTHESIZED_WIRE_749;
wire	SYNTHESIZED_WIRE_750;
wire	SYNTHESIZED_WIRE_751;
wire	SYNTHESIZED_WIRE_752;
wire	SYNTHESIZED_WIRE_753;
wire	SYNTHESIZED_WIRE_754;
wire	SYNTHESIZED_WIRE_755;
wire	SYNTHESIZED_WIRE_756;
wire	SYNTHESIZED_WIRE_757;
wire	SYNTHESIZED_WIRE_758;
wire	SYNTHESIZED_WIRE_759;
wire	SYNTHESIZED_WIRE_760;
wire	SYNTHESIZED_WIRE_761;
wire	SYNTHESIZED_WIRE_762;
wire	SYNTHESIZED_WIRE_763;
wire	SYNTHESIZED_WIRE_764;
wire	SYNTHESIZED_WIRE_765;
wire	SYNTHESIZED_WIRE_766;
wire	SYNTHESIZED_WIRE_767;
wire	SYNTHESIZED_WIRE_768;
wire	SYNTHESIZED_WIRE_769;
wire	SYNTHESIZED_WIRE_770;
wire	SYNTHESIZED_WIRE_771;
wire	SYNTHESIZED_WIRE_772;
wire	SYNTHESIZED_WIRE_773;
wire	SYNTHESIZED_WIRE_774;
wire	SYNTHESIZED_WIRE_775;
wire	SYNTHESIZED_WIRE_776;
wire	SYNTHESIZED_WIRE_777;
wire	SYNTHESIZED_WIRE_778;
wire	SYNTHESIZED_WIRE_779;
wire	SYNTHESIZED_WIRE_780;
wire	SYNTHESIZED_WIRE_781;
wire	SYNTHESIZED_WIRE_782;
wire	SYNTHESIZED_WIRE_783;
wire	SYNTHESIZED_WIRE_784;
wire	SYNTHESIZED_WIRE_785;
wire	SYNTHESIZED_WIRE_786;
wire	SYNTHESIZED_WIRE_787;
wire	SYNTHESIZED_WIRE_788;
wire	SYNTHESIZED_WIRE_789;
wire	SYNTHESIZED_WIRE_790;
wire	SYNTHESIZED_WIRE_791;
wire	SYNTHESIZED_WIRE_792;
wire	SYNTHESIZED_WIRE_793;
wire	SYNTHESIZED_WIRE_794;
wire	SYNTHESIZED_WIRE_795;
wire	SYNTHESIZED_WIRE_796;
wire	SYNTHESIZED_WIRE_797;
wire	SYNTHESIZED_WIRE_798;
wire	SYNTHESIZED_WIRE_799;
wire	SYNTHESIZED_WIRE_800;
wire	SYNTHESIZED_WIRE_801;
wire	SYNTHESIZED_WIRE_802;
wire	SYNTHESIZED_WIRE_803;
wire	SYNTHESIZED_WIRE_804;
wire	SYNTHESIZED_WIRE_805;
wire	SYNTHESIZED_WIRE_806;
wire	SYNTHESIZED_WIRE_807;
wire	SYNTHESIZED_WIRE_808;
wire	SYNTHESIZED_WIRE_809;
wire	SYNTHESIZED_WIRE_810;
wire	SYNTHESIZED_WIRE_811;
wire	SYNTHESIZED_WIRE_812;
wire	SYNTHESIZED_WIRE_813;
wire	SYNTHESIZED_WIRE_814;
wire	SYNTHESIZED_WIRE_815;
wire	SYNTHESIZED_WIRE_816;
wire	SYNTHESIZED_WIRE_817;
wire	SYNTHESIZED_WIRE_818;
wire	SYNTHESIZED_WIRE_819;
wire	SYNTHESIZED_WIRE_820;
wire	SYNTHESIZED_WIRE_821;
wire	SYNTHESIZED_WIRE_822;
wire	SYNTHESIZED_WIRE_823;
wire	SYNTHESIZED_WIRE_824;
wire	SYNTHESIZED_WIRE_825;
wire	SYNTHESIZED_WIRE_826;
wire	SYNTHESIZED_WIRE_827;
wire	SYNTHESIZED_WIRE_828;
wire	SYNTHESIZED_WIRE_829;
wire	SYNTHESIZED_WIRE_830;
wire	SYNTHESIZED_WIRE_831;
wire	SYNTHESIZED_WIRE_832;
wire	SYNTHESIZED_WIRE_833;
wire	SYNTHESIZED_WIRE_834;
wire	SYNTHESIZED_WIRE_835;
wire	SYNTHESIZED_WIRE_836;
wire	SYNTHESIZED_WIRE_837;
wire	SYNTHESIZED_WIRE_838;
wire	SYNTHESIZED_WIRE_839;
wire	SYNTHESIZED_WIRE_840;
wire	SYNTHESIZED_WIRE_841;
wire	SYNTHESIZED_WIRE_842;
wire	SYNTHESIZED_WIRE_843;
wire	SYNTHESIZED_WIRE_844;
wire	SYNTHESIZED_WIRE_845;
wire	SYNTHESIZED_WIRE_846;
wire	SYNTHESIZED_WIRE_847;
wire	SYNTHESIZED_WIRE_848;
wire	SYNTHESIZED_WIRE_849;
wire	SYNTHESIZED_WIRE_850;
wire	SYNTHESIZED_WIRE_851;
wire	SYNTHESIZED_WIRE_852;
wire	SYNTHESIZED_WIRE_853;
wire	SYNTHESIZED_WIRE_854;
wire	SYNTHESIZED_WIRE_855;
wire	SYNTHESIZED_WIRE_856;
wire	SYNTHESIZED_WIRE_857;
wire	SYNTHESIZED_WIRE_858;
wire	SYNTHESIZED_WIRE_859;
wire	SYNTHESIZED_WIRE_860;
wire	SYNTHESIZED_WIRE_861;
wire	SYNTHESIZED_WIRE_862;
wire	SYNTHESIZED_WIRE_863;
wire	SYNTHESIZED_WIRE_864;
wire	SYNTHESIZED_WIRE_865;
wire	SYNTHESIZED_WIRE_866;
wire	SYNTHESIZED_WIRE_867;
wire	SYNTHESIZED_WIRE_868;
wire	SYNTHESIZED_WIRE_869;
wire	SYNTHESIZED_WIRE_870;
wire	SYNTHESIZED_WIRE_871;
wire	SYNTHESIZED_WIRE_872;
wire	SYNTHESIZED_WIRE_873;
wire	SYNTHESIZED_WIRE_874;
wire	SYNTHESIZED_WIRE_875;
wire	SYNTHESIZED_WIRE_876;
wire	SYNTHESIZED_WIRE_877;
wire	SYNTHESIZED_WIRE_878;
wire	SYNTHESIZED_WIRE_879;
wire	SYNTHESIZED_WIRE_880;
wire	SYNTHESIZED_WIRE_881;
wire	SYNTHESIZED_WIRE_882;
wire	SYNTHESIZED_WIRE_883;
wire	SYNTHESIZED_WIRE_884;
wire	SYNTHESIZED_WIRE_885;
wire	SYNTHESIZED_WIRE_886;
wire	SYNTHESIZED_WIRE_887;
wire	SYNTHESIZED_WIRE_888;
wire	SYNTHESIZED_WIRE_889;
wire	SYNTHESIZED_WIRE_890;
wire	SYNTHESIZED_WIRE_891;
wire	SYNTHESIZED_WIRE_892;
wire	SYNTHESIZED_WIRE_893;
wire	SYNTHESIZED_WIRE_894;
wire	SYNTHESIZED_WIRE_895;
wire	SYNTHESIZED_WIRE_896;
wire	SYNTHESIZED_WIRE_897;
wire	SYNTHESIZED_WIRE_898;
wire	SYNTHESIZED_WIRE_899;
wire	SYNTHESIZED_WIRE_900;
wire	SYNTHESIZED_WIRE_901;
wire	SYNTHESIZED_WIRE_902;
wire	SYNTHESIZED_WIRE_903;
wire	SYNTHESIZED_WIRE_904;
wire	SYNTHESIZED_WIRE_905;
wire	SYNTHESIZED_WIRE_906;
wire	SYNTHESIZED_WIRE_907;
wire	SYNTHESIZED_WIRE_908;
wire	SYNTHESIZED_WIRE_909;
wire	SYNTHESIZED_WIRE_910;
wire	SYNTHESIZED_WIRE_911;
wire	SYNTHESIZED_WIRE_912;
wire	SYNTHESIZED_WIRE_913;
wire	SYNTHESIZED_WIRE_914;
wire	SYNTHESIZED_WIRE_915;
wire	SYNTHESIZED_WIRE_916;
wire	SYNTHESIZED_WIRE_917;
wire	SYNTHESIZED_WIRE_918;
wire	SYNTHESIZED_WIRE_919;
wire	SYNTHESIZED_WIRE_920;
wire	SYNTHESIZED_WIRE_921;
wire	SYNTHESIZED_WIRE_922;
wire	SYNTHESIZED_WIRE_923;
wire	SYNTHESIZED_WIRE_924;
wire	SYNTHESIZED_WIRE_925;
wire	SYNTHESIZED_WIRE_926;
wire	SYNTHESIZED_WIRE_927;
wire	SYNTHESIZED_WIRE_928;
wire	SYNTHESIZED_WIRE_929;
wire	SYNTHESIZED_WIRE_930;
wire	SYNTHESIZED_WIRE_931;
wire	SYNTHESIZED_WIRE_932;
wire	SYNTHESIZED_WIRE_933;
wire	SYNTHESIZED_WIRE_934;
wire	SYNTHESIZED_WIRE_935;
wire	SYNTHESIZED_WIRE_936;
wire	SYNTHESIZED_WIRE_937;
wire	SYNTHESIZED_WIRE_938;
wire	SYNTHESIZED_WIRE_939;
wire	SYNTHESIZED_WIRE_940;
wire	SYNTHESIZED_WIRE_941;
wire	SYNTHESIZED_WIRE_942;
wire	SYNTHESIZED_WIRE_943;
wire	SYNTHESIZED_WIRE_944;
wire	SYNTHESIZED_WIRE_945;
wire	SYNTHESIZED_WIRE_946;
wire	SYNTHESIZED_WIRE_947;
wire	SYNTHESIZED_WIRE_948;
wire	SYNTHESIZED_WIRE_949;
wire	SYNTHESIZED_WIRE_950;
wire	SYNTHESIZED_WIRE_951;
wire	SYNTHESIZED_WIRE_952;
wire	SYNTHESIZED_WIRE_953;
wire	SYNTHESIZED_WIRE_954;
wire	SYNTHESIZED_WIRE_955;
wire	SYNTHESIZED_WIRE_956;
wire	SYNTHESIZED_WIRE_957;
wire	SYNTHESIZED_WIRE_958;
wire	SYNTHESIZED_WIRE_959;
wire	SYNTHESIZED_WIRE_960;
wire	SYNTHESIZED_WIRE_961;
wire	SYNTHESIZED_WIRE_962;
wire	SYNTHESIZED_WIRE_963;
wire	SYNTHESIZED_WIRE_964;
wire	SYNTHESIZED_WIRE_965;
wire	SYNTHESIZED_WIRE_966;
wire	SYNTHESIZED_WIRE_967;
wire	SYNTHESIZED_WIRE_968;
wire	SYNTHESIZED_WIRE_969;
wire	SYNTHESIZED_WIRE_970;
wire	SYNTHESIZED_WIRE_971;
wire	SYNTHESIZED_WIRE_972;
wire	SYNTHESIZED_WIRE_973;
wire	SYNTHESIZED_WIRE_974;
wire	SYNTHESIZED_WIRE_975;
wire	SYNTHESIZED_WIRE_976;
wire	SYNTHESIZED_WIRE_977;
wire	SYNTHESIZED_WIRE_978;
wire	SYNTHESIZED_WIRE_979;
wire	SYNTHESIZED_WIRE_980;
wire	SYNTHESIZED_WIRE_981;
wire	SYNTHESIZED_WIRE_982;
wire	SYNTHESIZED_WIRE_983;
wire	SYNTHESIZED_WIRE_984;
wire	SYNTHESIZED_WIRE_985;
wire	SYNTHESIZED_WIRE_986;
wire	SYNTHESIZED_WIRE_987;
wire	SYNTHESIZED_WIRE_988;
wire	SYNTHESIZED_WIRE_989;
wire	SYNTHESIZED_WIRE_990;
wire	SYNTHESIZED_WIRE_991;
wire	SYNTHESIZED_WIRE_992;
wire	SYNTHESIZED_WIRE_993;
wire	SYNTHESIZED_WIRE_994;
wire	SYNTHESIZED_WIRE_995;
wire	SYNTHESIZED_WIRE_996;
wire	SYNTHESIZED_WIRE_997;
wire	SYNTHESIZED_WIRE_998;
wire	SYNTHESIZED_WIRE_999;
wire	SYNTHESIZED_WIRE_1000;
wire	SYNTHESIZED_WIRE_1001;
wire	SYNTHESIZED_WIRE_1002;
wire	SYNTHESIZED_WIRE_1003;
wire	SYNTHESIZED_WIRE_1004;
wire	SYNTHESIZED_WIRE_1005;
wire	SYNTHESIZED_WIRE_1006;
wire	SYNTHESIZED_WIRE_1007;
wire	SYNTHESIZED_WIRE_1008;
wire	SYNTHESIZED_WIRE_1009;
wire	SYNTHESIZED_WIRE_1010;
wire	SYNTHESIZED_WIRE_1011;
wire	SYNTHESIZED_WIRE_1012;
wire	SYNTHESIZED_WIRE_1013;
wire	SYNTHESIZED_WIRE_1014;
wire	SYNTHESIZED_WIRE_1015;
wire	SYNTHESIZED_WIRE_1016;
wire	SYNTHESIZED_WIRE_1017;
wire	SYNTHESIZED_WIRE_1018;
wire	SYNTHESIZED_WIRE_1019;
wire	SYNTHESIZED_WIRE_1020;
wire	SYNTHESIZED_WIRE_1021;
wire	SYNTHESIZED_WIRE_1022;
wire	SYNTHESIZED_WIRE_1023;
wire	SYNTHESIZED_WIRE_1024;
wire	SYNTHESIZED_WIRE_1025;
wire	SYNTHESIZED_WIRE_1026;
wire	SYNTHESIZED_WIRE_1027;
wire	SYNTHESIZED_WIRE_1028;
wire	SYNTHESIZED_WIRE_1029;
wire	SYNTHESIZED_WIRE_1030;
wire	SYNTHESIZED_WIRE_1031;
wire	SYNTHESIZED_WIRE_1032;
wire	SYNTHESIZED_WIRE_1033;
wire	SYNTHESIZED_WIRE_1034;
wire	SYNTHESIZED_WIRE_1035;
wire	SYNTHESIZED_WIRE_1036;
wire	SYNTHESIZED_WIRE_1037;
wire	SYNTHESIZED_WIRE_1038;
wire	SYNTHESIZED_WIRE_1039;
wire	SYNTHESIZED_WIRE_1040;
wire	SYNTHESIZED_WIRE_1041;
wire	SYNTHESIZED_WIRE_1042;
wire	SYNTHESIZED_WIRE_1043;
wire	SYNTHESIZED_WIRE_1044;
wire	SYNTHESIZED_WIRE_1045;
wire	SYNTHESIZED_WIRE_1046;
wire	SYNTHESIZED_WIRE_1047;
wire	SYNTHESIZED_WIRE_1048;
wire	SYNTHESIZED_WIRE_1049;
wire	SYNTHESIZED_WIRE_1050;
wire	SYNTHESIZED_WIRE_1051;
wire	SYNTHESIZED_WIRE_1052;
wire	SYNTHESIZED_WIRE_1053;
wire	SYNTHESIZED_WIRE_1054;
wire	SYNTHESIZED_WIRE_1055;
wire	SYNTHESIZED_WIRE_1056;
wire	SYNTHESIZED_WIRE_1057;
wire	SYNTHESIZED_WIRE_1058;
wire	SYNTHESIZED_WIRE_1059;
wire	SYNTHESIZED_WIRE_1060;
wire	SYNTHESIZED_WIRE_1061;
wire	SYNTHESIZED_WIRE_1062;
wire	SYNTHESIZED_WIRE_1063;
wire	SYNTHESIZED_WIRE_1064;
wire	SYNTHESIZED_WIRE_1065;
wire	SYNTHESIZED_WIRE_1066;
wire	SYNTHESIZED_WIRE_1067;
wire	SYNTHESIZED_WIRE_1068;
wire	SYNTHESIZED_WIRE_1069;
wire	SYNTHESIZED_WIRE_1070;
wire	SYNTHESIZED_WIRE_1071;
wire	SYNTHESIZED_WIRE_1072;
wire	SYNTHESIZED_WIRE_1073;
wire	SYNTHESIZED_WIRE_1074;
wire	SYNTHESIZED_WIRE_1075;
wire	SYNTHESIZED_WIRE_1076;
wire	SYNTHESIZED_WIRE_1077;
wire	SYNTHESIZED_WIRE_1078;
wire	SYNTHESIZED_WIRE_1079;
wire	SYNTHESIZED_WIRE_1080;
wire	SYNTHESIZED_WIRE_1081;
wire	SYNTHESIZED_WIRE_1082;
wire	SYNTHESIZED_WIRE_1083;
wire	SYNTHESIZED_WIRE_1084;
wire	SYNTHESIZED_WIRE_1085;
wire	SYNTHESIZED_WIRE_1086;
wire	SYNTHESIZED_WIRE_1087;
wire	SYNTHESIZED_WIRE_1088;
wire	SYNTHESIZED_WIRE_1089;
wire	SYNTHESIZED_WIRE_1090;
wire	SYNTHESIZED_WIRE_1091;
wire	SYNTHESIZED_WIRE_1092;
wire	SYNTHESIZED_WIRE_1093;
wire	SYNTHESIZED_WIRE_1094;
wire	SYNTHESIZED_WIRE_1095;
wire	SYNTHESIZED_WIRE_1096;
wire	SYNTHESIZED_WIRE_1097;
wire	SYNTHESIZED_WIRE_1098;
wire	SYNTHESIZED_WIRE_1099;
wire	SYNTHESIZED_WIRE_1100;
wire	SYNTHESIZED_WIRE_1101;
wire	SYNTHESIZED_WIRE_1102;
wire	SYNTHESIZED_WIRE_1103;
wire	SYNTHESIZED_WIRE_1104;
wire	SYNTHESIZED_WIRE_1105;
wire	SYNTHESIZED_WIRE_1106;
wire	SYNTHESIZED_WIRE_1107;
wire	SYNTHESIZED_WIRE_1108;
wire	SYNTHESIZED_WIRE_1109;
wire	SYNTHESIZED_WIRE_1110;
wire	SYNTHESIZED_WIRE_1111;
wire	SYNTHESIZED_WIRE_1112;
wire	SYNTHESIZED_WIRE_1113;
wire	SYNTHESIZED_WIRE_1114;
wire	SYNTHESIZED_WIRE_1115;
wire	SYNTHESIZED_WIRE_1116;
wire	SYNTHESIZED_WIRE_1117;
wire	SYNTHESIZED_WIRE_1118;
wire	SYNTHESIZED_WIRE_1119;
wire	SYNTHESIZED_WIRE_1120;
wire	SYNTHESIZED_WIRE_1121;
wire	SYNTHESIZED_WIRE_1122;
wire	SYNTHESIZED_WIRE_1123;
wire	SYNTHESIZED_WIRE_1124;
wire	SYNTHESIZED_WIRE_1125;
wire	SYNTHESIZED_WIRE_1126;
wire	SYNTHESIZED_WIRE_1127;
wire	SYNTHESIZED_WIRE_1128;
wire	SYNTHESIZED_WIRE_1129;
wire	SYNTHESIZED_WIRE_1130;
wire	SYNTHESIZED_WIRE_1131;
wire	SYNTHESIZED_WIRE_1132;
wire	SYNTHESIZED_WIRE_1133;
wire	SYNTHESIZED_WIRE_1134;
wire	SYNTHESIZED_WIRE_1135;
wire	SYNTHESIZED_WIRE_1136;
wire	SYNTHESIZED_WIRE_1137;
wire	SYNTHESIZED_WIRE_1138;
wire	SYNTHESIZED_WIRE_1139;
wire	SYNTHESIZED_WIRE_1140;
wire	SYNTHESIZED_WIRE_1141;
wire	SYNTHESIZED_WIRE_1142;
wire	SYNTHESIZED_WIRE_1143;
wire	SYNTHESIZED_WIRE_1144;
wire	SYNTHESIZED_WIRE_1145;
wire	SYNTHESIZED_WIRE_1146;
wire	SYNTHESIZED_WIRE_1147;
wire	SYNTHESIZED_WIRE_1148;
wire	SYNTHESIZED_WIRE_1149;
wire	SYNTHESIZED_WIRE_1150;
wire	SYNTHESIZED_WIRE_1151;
wire	SYNTHESIZED_WIRE_1152;
wire	SYNTHESIZED_WIRE_1153;
wire	SYNTHESIZED_WIRE_1154;
wire	SYNTHESIZED_WIRE_1155;
wire	SYNTHESIZED_WIRE_1156;
wire	SYNTHESIZED_WIRE_1157;
wire	SYNTHESIZED_WIRE_1158;
wire	SYNTHESIZED_WIRE_1159;
wire	SYNTHESIZED_WIRE_1160;
wire	SYNTHESIZED_WIRE_1161;
wire	SYNTHESIZED_WIRE_1162;
wire	SYNTHESIZED_WIRE_1163;
wire	SYNTHESIZED_WIRE_1164;
wire	SYNTHESIZED_WIRE_1165;
wire	SYNTHESIZED_WIRE_1166;
wire	SYNTHESIZED_WIRE_1167;
wire	SYNTHESIZED_WIRE_1168;
wire	SYNTHESIZED_WIRE_1169;
wire	SYNTHESIZED_WIRE_1170;
wire	SYNTHESIZED_WIRE_1171;
wire	SYNTHESIZED_WIRE_1172;
wire	SYNTHESIZED_WIRE_1173;
wire	SYNTHESIZED_WIRE_1174;
wire	SYNTHESIZED_WIRE_1175;
wire	SYNTHESIZED_WIRE_1176;
wire	SYNTHESIZED_WIRE_1177;
wire	SYNTHESIZED_WIRE_1178;
wire	SYNTHESIZED_WIRE_1179;
wire	SYNTHESIZED_WIRE_1180;
wire	SYNTHESIZED_WIRE_1181;
wire	SYNTHESIZED_WIRE_1182;
wire	SYNTHESIZED_WIRE_1183;
wire	SYNTHESIZED_WIRE_1184;
wire	SYNTHESIZED_WIRE_1185;
wire	SYNTHESIZED_WIRE_1186;
wire	SYNTHESIZED_WIRE_1187;
wire	SYNTHESIZED_WIRE_1188;
wire	SYNTHESIZED_WIRE_1189;
wire	SYNTHESIZED_WIRE_1190;
wire	SYNTHESIZED_WIRE_1191;
wire	SYNTHESIZED_WIRE_1192;
wire	SYNTHESIZED_WIRE_1193;
wire	SYNTHESIZED_WIRE_1194;
wire	SYNTHESIZED_WIRE_1195;
wire	SYNTHESIZED_WIRE_1196;
wire	SYNTHESIZED_WIRE_1197;
wire	SYNTHESIZED_WIRE_1198;
wire	SYNTHESIZED_WIRE_1199;
wire	SYNTHESIZED_WIRE_1200;
wire	SYNTHESIZED_WIRE_1201;
wire	SYNTHESIZED_WIRE_1202;
wire	SYNTHESIZED_WIRE_1203;
wire	SYNTHESIZED_WIRE_1204;
wire	SYNTHESIZED_WIRE_1205;
wire	SYNTHESIZED_WIRE_1206;
wire	SYNTHESIZED_WIRE_1207;
wire	SYNTHESIZED_WIRE_1208;
wire	SYNTHESIZED_WIRE_1209;
wire	SYNTHESIZED_WIRE_1210;
wire	SYNTHESIZED_WIRE_1211;
wire	SYNTHESIZED_WIRE_1212;
wire	SYNTHESIZED_WIRE_1213;
wire	SYNTHESIZED_WIRE_1214;
wire	SYNTHESIZED_WIRE_1215;
wire	SYNTHESIZED_WIRE_1216;
wire	SYNTHESIZED_WIRE_1217;
wire	SYNTHESIZED_WIRE_1218;
wire	SYNTHESIZED_WIRE_1219;
wire	SYNTHESIZED_WIRE_1220;
wire	SYNTHESIZED_WIRE_1221;
wire	SYNTHESIZED_WIRE_1222;
wire	SYNTHESIZED_WIRE_1223;
wire	SYNTHESIZED_WIRE_1224;
wire	SYNTHESIZED_WIRE_1225;
wire	SYNTHESIZED_WIRE_1226;
wire	SYNTHESIZED_WIRE_1227;
wire	SYNTHESIZED_WIRE_1228;
wire	SYNTHESIZED_WIRE_1229;
wire	SYNTHESIZED_WIRE_1230;
wire	SYNTHESIZED_WIRE_1231;
wire	SYNTHESIZED_WIRE_1232;
wire	SYNTHESIZED_WIRE_1233;
wire	SYNTHESIZED_WIRE_1234;
wire	SYNTHESIZED_WIRE_1235;
wire	SYNTHESIZED_WIRE_1236;
wire	SYNTHESIZED_WIRE_1237;
wire	SYNTHESIZED_WIRE_1238;
wire	SYNTHESIZED_WIRE_1239;
wire	SYNTHESIZED_WIRE_1240;
wire	SYNTHESIZED_WIRE_1241;
wire	SYNTHESIZED_WIRE_1242;
wire	SYNTHESIZED_WIRE_1243;
wire	SYNTHESIZED_WIRE_1244;
wire	SYNTHESIZED_WIRE_1245;
wire	SYNTHESIZED_WIRE_1246;
wire	SYNTHESIZED_WIRE_1247;
wire	SYNTHESIZED_WIRE_1248;
wire	SYNTHESIZED_WIRE_1249;
wire	SYNTHESIZED_WIRE_1250;
wire	SYNTHESIZED_WIRE_1251;
wire	SYNTHESIZED_WIRE_1252;
wire	SYNTHESIZED_WIRE_1253;
wire	SYNTHESIZED_WIRE_1254;
wire	SYNTHESIZED_WIRE_1255;
wire	SYNTHESIZED_WIRE_1256;
wire	SYNTHESIZED_WIRE_1257;
wire	SYNTHESIZED_WIRE_1258;
wire	SYNTHESIZED_WIRE_1259;
wire	SYNTHESIZED_WIRE_1260;
wire	SYNTHESIZED_WIRE_1261;
wire	SYNTHESIZED_WIRE_1262;
wire	SYNTHESIZED_WIRE_1263;
wire	SYNTHESIZED_WIRE_1264;
wire	SYNTHESIZED_WIRE_1265;
wire	SYNTHESIZED_WIRE_1266;
wire	SYNTHESIZED_WIRE_1267;
wire	SYNTHESIZED_WIRE_1268;
wire	SYNTHESIZED_WIRE_1269;
wire	SYNTHESIZED_WIRE_1270;
wire	SYNTHESIZED_WIRE_1271;
wire	SYNTHESIZED_WIRE_1272;
wire	SYNTHESIZED_WIRE_1273;
wire	SYNTHESIZED_WIRE_1274;
wire	SYNTHESIZED_WIRE_1275;
wire	SYNTHESIZED_WIRE_1276;
wire	SYNTHESIZED_WIRE_1277;
wire	SYNTHESIZED_WIRE_1278;
wire	SYNTHESIZED_WIRE_1279;
wire	SYNTHESIZED_WIRE_1280;
wire	SYNTHESIZED_WIRE_1281;
wire	SYNTHESIZED_WIRE_1282;
wire	SYNTHESIZED_WIRE_1283;
wire	SYNTHESIZED_WIRE_1284;
wire	SYNTHESIZED_WIRE_1285;
wire	SYNTHESIZED_WIRE_1286;
wire	SYNTHESIZED_WIRE_1287;
wire	SYNTHESIZED_WIRE_1288;
wire	SYNTHESIZED_WIRE_1289;
wire	SYNTHESIZED_WIRE_1290;
wire	SYNTHESIZED_WIRE_1291;
wire	SYNTHESIZED_WIRE_1292;
wire	SYNTHESIZED_WIRE_1293;
wire	SYNTHESIZED_WIRE_1294;
wire	SYNTHESIZED_WIRE_1295;
wire	SYNTHESIZED_WIRE_1296;
wire	SYNTHESIZED_WIRE_1297;
wire	SYNTHESIZED_WIRE_1298;
wire	SYNTHESIZED_WIRE_1299;
wire	SYNTHESIZED_WIRE_1300;
wire	SYNTHESIZED_WIRE_1301;
wire	SYNTHESIZED_WIRE_1302;
wire	SYNTHESIZED_WIRE_1303;
wire	SYNTHESIZED_WIRE_1304;
wire	SYNTHESIZED_WIRE_1305;
wire	SYNTHESIZED_WIRE_1306;
wire	SYNTHESIZED_WIRE_1307;
wire	SYNTHESIZED_WIRE_1308;
wire	SYNTHESIZED_WIRE_1309;
wire	SYNTHESIZED_WIRE_1310;
wire	SYNTHESIZED_WIRE_1311;
wire	SYNTHESIZED_WIRE_1312;
wire	SYNTHESIZED_WIRE_1313;
wire	SYNTHESIZED_WIRE_1314;
wire	SYNTHESIZED_WIRE_1315;
wire	SYNTHESIZED_WIRE_1316;
wire	SYNTHESIZED_WIRE_1317;
wire	SYNTHESIZED_WIRE_1318;
wire	SYNTHESIZED_WIRE_1319;
wire	SYNTHESIZED_WIRE_1320;
wire	SYNTHESIZED_WIRE_1321;
wire	SYNTHESIZED_WIRE_1322;
wire	SYNTHESIZED_WIRE_1323;
wire	SYNTHESIZED_WIRE_1324;
wire	SYNTHESIZED_WIRE_1325;
wire	SYNTHESIZED_WIRE_1326;
wire	SYNTHESIZED_WIRE_1327;
wire	SYNTHESIZED_WIRE_1328;
wire	SYNTHESIZED_WIRE_1329;
wire	SYNTHESIZED_WIRE_1330;
wire	SYNTHESIZED_WIRE_1331;
wire	SYNTHESIZED_WIRE_1332;
wire	SYNTHESIZED_WIRE_1333;
wire	SYNTHESIZED_WIRE_1334;
wire	SYNTHESIZED_WIRE_1335;
wire	SYNTHESIZED_WIRE_1336;
wire	SYNTHESIZED_WIRE_1337;
wire	SYNTHESIZED_WIRE_1338;
wire	SYNTHESIZED_WIRE_1339;
wire	SYNTHESIZED_WIRE_1340;
wire	SYNTHESIZED_WIRE_1341;
wire	SYNTHESIZED_WIRE_1342;
wire	SYNTHESIZED_WIRE_1343;
wire	SYNTHESIZED_WIRE_1344;
wire	SYNTHESIZED_WIRE_1345;
wire	SYNTHESIZED_WIRE_1346;
wire	SYNTHESIZED_WIRE_1347;
wire	SYNTHESIZED_WIRE_1348;
wire	SYNTHESIZED_WIRE_1349;
wire	SYNTHESIZED_WIRE_1350;
wire	SYNTHESIZED_WIRE_1351;
wire	SYNTHESIZED_WIRE_1352;
wire	SYNTHESIZED_WIRE_1353;
wire	SYNTHESIZED_WIRE_1354;
wire	SYNTHESIZED_WIRE_1355;
wire	SYNTHESIZED_WIRE_1356;
wire	SYNTHESIZED_WIRE_1357;
wire	SYNTHESIZED_WIRE_1358;
wire	SYNTHESIZED_WIRE_1359;
wire	SYNTHESIZED_WIRE_1360;
wire	SYNTHESIZED_WIRE_1361;
wire	SYNTHESIZED_WIRE_1362;
wire	SYNTHESIZED_WIRE_1363;
wire	SYNTHESIZED_WIRE_1364;
wire	SYNTHESIZED_WIRE_1365;
wire	SYNTHESIZED_WIRE_1366;
wire	SYNTHESIZED_WIRE_1367;
wire	SYNTHESIZED_WIRE_1368;
wire	SYNTHESIZED_WIRE_1369;
wire	SYNTHESIZED_WIRE_1370;
wire	SYNTHESIZED_WIRE_1371;
wire	SYNTHESIZED_WIRE_1372;
wire	SYNTHESIZED_WIRE_1373;
wire	SYNTHESIZED_WIRE_1374;
wire	SYNTHESIZED_WIRE_1375;
wire	SYNTHESIZED_WIRE_1376;
wire	SYNTHESIZED_WIRE_1377;
wire	SYNTHESIZED_WIRE_1378;
wire	SYNTHESIZED_WIRE_1379;
wire	SYNTHESIZED_WIRE_1380;
wire	SYNTHESIZED_WIRE_1381;
wire	SYNTHESIZED_WIRE_1382;
wire	SYNTHESIZED_WIRE_1383;
wire	SYNTHESIZED_WIRE_1384;
wire	SYNTHESIZED_WIRE_1385;
wire	SYNTHESIZED_WIRE_1386;
wire	SYNTHESIZED_WIRE_1387;
wire	SYNTHESIZED_WIRE_1388;
wire	SYNTHESIZED_WIRE_1389;
wire	SYNTHESIZED_WIRE_1390;
wire	SYNTHESIZED_WIRE_1391;
wire	SYNTHESIZED_WIRE_1392;
wire	SYNTHESIZED_WIRE_1393;
wire	SYNTHESIZED_WIRE_1394;
wire	SYNTHESIZED_WIRE_1395;
wire	SYNTHESIZED_WIRE_1396;
wire	SYNTHESIZED_WIRE_1397;
wire	SYNTHESIZED_WIRE_1398;
wire	SYNTHESIZED_WIRE_1399;
wire	SYNTHESIZED_WIRE_1400;
wire	SYNTHESIZED_WIRE_1401;
wire	SYNTHESIZED_WIRE_1402;
wire	SYNTHESIZED_WIRE_1403;
wire	SYNTHESIZED_WIRE_1404;
wire	SYNTHESIZED_WIRE_1405;
wire	SYNTHESIZED_WIRE_1406;
wire	SYNTHESIZED_WIRE_1407;
wire	SYNTHESIZED_WIRE_1408;
wire	SYNTHESIZED_WIRE_1409;
wire	SYNTHESIZED_WIRE_1410;
wire	SYNTHESIZED_WIRE_1411;
wire	SYNTHESIZED_WIRE_1412;
wire	SYNTHESIZED_WIRE_1413;
wire	SYNTHESIZED_WIRE_1414;
wire	SYNTHESIZED_WIRE_1415;
wire	SYNTHESIZED_WIRE_1416;
wire	SYNTHESIZED_WIRE_1417;
wire	SYNTHESIZED_WIRE_1418;
wire	SYNTHESIZED_WIRE_1419;
wire	SYNTHESIZED_WIRE_1420;
wire	SYNTHESIZED_WIRE_1421;
wire	SYNTHESIZED_WIRE_1422;
wire	SYNTHESIZED_WIRE_1423;
wire	SYNTHESIZED_WIRE_1424;
wire	SYNTHESIZED_WIRE_1425;
wire	SYNTHESIZED_WIRE_1426;
wire	SYNTHESIZED_WIRE_1427;
wire	SYNTHESIZED_WIRE_1428;
wire	SYNTHESIZED_WIRE_1429;
wire	SYNTHESIZED_WIRE_1430;
wire	SYNTHESIZED_WIRE_1431;
wire	SYNTHESIZED_WIRE_1432;
wire	SYNTHESIZED_WIRE_1433;
wire	SYNTHESIZED_WIRE_1434;
wire	SYNTHESIZED_WIRE_1435;
wire	SYNTHESIZED_WIRE_1436;
wire	SYNTHESIZED_WIRE_1437;
wire	SYNTHESIZED_WIRE_1438;
wire	SYNTHESIZED_WIRE_1439;
wire	SYNTHESIZED_WIRE_1440;
wire	SYNTHESIZED_WIRE_1441;
wire	SYNTHESIZED_WIRE_1442;
wire	SYNTHESIZED_WIRE_1443;
wire	SYNTHESIZED_WIRE_1444;
wire	SYNTHESIZED_WIRE_1445;
wire	SYNTHESIZED_WIRE_1446;
wire	SYNTHESIZED_WIRE_1447;
wire	SYNTHESIZED_WIRE_1448;
wire	SYNTHESIZED_WIRE_1449;
wire	SYNTHESIZED_WIRE_1450;
wire	SYNTHESIZED_WIRE_1451;
wire	SYNTHESIZED_WIRE_1452;
wire	SYNTHESIZED_WIRE_1453;
wire	SYNTHESIZED_WIRE_1454;
wire	SYNTHESIZED_WIRE_1455;
wire	SYNTHESIZED_WIRE_1456;
wire	SYNTHESIZED_WIRE_1457;
wire	SYNTHESIZED_WIRE_1458;
wire	SYNTHESIZED_WIRE_1459;
wire	SYNTHESIZED_WIRE_1460;
wire	SYNTHESIZED_WIRE_1461;
wire	SYNTHESIZED_WIRE_1462;
wire	SYNTHESIZED_WIRE_1463;
wire	SYNTHESIZED_WIRE_1464;
wire	SYNTHESIZED_WIRE_1465;
wire	SYNTHESIZED_WIRE_1466;
wire	SYNTHESIZED_WIRE_1467;
wire	SYNTHESIZED_WIRE_1468;
wire	SYNTHESIZED_WIRE_1469;
wire	SYNTHESIZED_WIRE_1470;
wire	SYNTHESIZED_WIRE_1471;
wire	SYNTHESIZED_WIRE_1472;
wire	SYNTHESIZED_WIRE_1473;
wire	SYNTHESIZED_WIRE_1474;
wire	SYNTHESIZED_WIRE_1475;
wire	SYNTHESIZED_WIRE_1476;
wire	SYNTHESIZED_WIRE_1477;
wire	SYNTHESIZED_WIRE_1478;
wire	SYNTHESIZED_WIRE_1479;
wire	SYNTHESIZED_WIRE_1480;
wire	SYNTHESIZED_WIRE_1481;
wire	SYNTHESIZED_WIRE_1482;
wire	SYNTHESIZED_WIRE_1483;
wire	SYNTHESIZED_WIRE_1484;
wire	SYNTHESIZED_WIRE_1485;
wire	SYNTHESIZED_WIRE_1486;
wire	SYNTHESIZED_WIRE_1487;
wire	SYNTHESIZED_WIRE_1488;
wire	SYNTHESIZED_WIRE_1489;
wire	SYNTHESIZED_WIRE_1490;
wire	SYNTHESIZED_WIRE_1491;
wire	SYNTHESIZED_WIRE_1492;
wire	SYNTHESIZED_WIRE_1493;
wire	SYNTHESIZED_WIRE_1494;
wire	SYNTHESIZED_WIRE_1495;
wire	SYNTHESIZED_WIRE_1496;
wire	SYNTHESIZED_WIRE_1497;
wire	SYNTHESIZED_WIRE_1498;
wire	SYNTHESIZED_WIRE_1499;
wire	SYNTHESIZED_WIRE_1500;
wire	SYNTHESIZED_WIRE_1501;
wire	SYNTHESIZED_WIRE_1502;
wire	SYNTHESIZED_WIRE_1503;
wire	SYNTHESIZED_WIRE_1504;
wire	SYNTHESIZED_WIRE_1505;
wire	SYNTHESIZED_WIRE_1506;
wire	SYNTHESIZED_WIRE_1507;
wire	SYNTHESIZED_WIRE_1508;
wire	SYNTHESIZED_WIRE_1509;
wire	SYNTHESIZED_WIRE_1510;
wire	SYNTHESIZED_WIRE_1511;
wire	SYNTHESIZED_WIRE_1512;
wire	SYNTHESIZED_WIRE_1513;
wire	SYNTHESIZED_WIRE_1514;
wire	SYNTHESIZED_WIRE_1515;
wire	SYNTHESIZED_WIRE_1516;
wire	SYNTHESIZED_WIRE_1517;
wire	SYNTHESIZED_WIRE_1518;
wire	SYNTHESIZED_WIRE_1519;
wire	SYNTHESIZED_WIRE_1520;
wire	SYNTHESIZED_WIRE_1521;
wire	SYNTHESIZED_WIRE_1522;
wire	SYNTHESIZED_WIRE_1523;
wire	SYNTHESIZED_WIRE_1524;
wire	SYNTHESIZED_WIRE_1525;
wire	SYNTHESIZED_WIRE_1526;
wire	SYNTHESIZED_WIRE_1527;
wire	SYNTHESIZED_WIRE_1528;
wire	SYNTHESIZED_WIRE_1529;
wire	SYNTHESIZED_WIRE_1530;
wire	SYNTHESIZED_WIRE_1531;
wire	SYNTHESIZED_WIRE_1532;
wire	SYNTHESIZED_WIRE_1533;
wire	SYNTHESIZED_WIRE_1534;
wire	SYNTHESIZED_WIRE_1535;
wire	SYNTHESIZED_WIRE_1536;
wire	SYNTHESIZED_WIRE_1537;
wire	SYNTHESIZED_WIRE_1538;
wire	SYNTHESIZED_WIRE_1539;
wire	SYNTHESIZED_WIRE_1540;
wire	SYNTHESIZED_WIRE_1541;
wire	SYNTHESIZED_WIRE_1542;
wire	SYNTHESIZED_WIRE_1543;
wire	SYNTHESIZED_WIRE_1544;
wire	SYNTHESIZED_WIRE_1545;
wire	SYNTHESIZED_WIRE_1546;
wire	SYNTHESIZED_WIRE_1547;
wire	SYNTHESIZED_WIRE_1548;
wire	SYNTHESIZED_WIRE_1549;
wire	SYNTHESIZED_WIRE_1550;
wire	SYNTHESIZED_WIRE_1551;
wire	SYNTHESIZED_WIRE_1552;
wire	SYNTHESIZED_WIRE_1553;
wire	SYNTHESIZED_WIRE_1554;
wire	SYNTHESIZED_WIRE_1555;
wire	SYNTHESIZED_WIRE_1556;
wire	SYNTHESIZED_WIRE_1557;
wire	SYNTHESIZED_WIRE_1558;
wire	SYNTHESIZED_WIRE_1559;
wire	SYNTHESIZED_WIRE_1560;
wire	SYNTHESIZED_WIRE_1561;
wire	SYNTHESIZED_WIRE_1562;
wire	SYNTHESIZED_WIRE_1563;
wire	SYNTHESIZED_WIRE_1564;
wire	SYNTHESIZED_WIRE_1565;
wire	SYNTHESIZED_WIRE_1566;
wire	SYNTHESIZED_WIRE_1567;
wire	SYNTHESIZED_WIRE_1568;
wire	SYNTHESIZED_WIRE_1569;
wire	SYNTHESIZED_WIRE_1570;
wire	SYNTHESIZED_WIRE_1571;
wire	SYNTHESIZED_WIRE_1572;
wire	SYNTHESIZED_WIRE_1573;
wire	SYNTHESIZED_WIRE_1574;
wire	SYNTHESIZED_WIRE_1575;
wire	SYNTHESIZED_WIRE_1576;
wire	SYNTHESIZED_WIRE_1577;
wire	SYNTHESIZED_WIRE_1578;
wire	SYNTHESIZED_WIRE_1579;
wire	SYNTHESIZED_WIRE_1580;
wire	SYNTHESIZED_WIRE_1581;
wire	SYNTHESIZED_WIRE_1582;
wire	SYNTHESIZED_WIRE_1583;
wire	SYNTHESIZED_WIRE_1584;
wire	SYNTHESIZED_WIRE_1585;
wire	SYNTHESIZED_WIRE_1586;
wire	SYNTHESIZED_WIRE_1587;
wire	SYNTHESIZED_WIRE_1588;
wire	SYNTHESIZED_WIRE_1589;
wire	SYNTHESIZED_WIRE_1590;
wire	SYNTHESIZED_WIRE_1591;
wire	SYNTHESIZED_WIRE_1592;
wire	SYNTHESIZED_WIRE_1593;
wire	SYNTHESIZED_WIRE_1594;
wire	SYNTHESIZED_WIRE_1595;
wire	SYNTHESIZED_WIRE_1596;
wire	SYNTHESIZED_WIRE_1597;
wire	SYNTHESIZED_WIRE_1598;
wire	SYNTHESIZED_WIRE_1599;
wire	SYNTHESIZED_WIRE_1600;
wire	SYNTHESIZED_WIRE_1601;
wire	SYNTHESIZED_WIRE_1602;
wire	SYNTHESIZED_WIRE_1603;
wire	SYNTHESIZED_WIRE_1604;
wire	SYNTHESIZED_WIRE_1605;
wire	SYNTHESIZED_WIRE_1606;
wire	SYNTHESIZED_WIRE_1607;
wire	SYNTHESIZED_WIRE_1608;
wire	SYNTHESIZED_WIRE_1609;
wire	SYNTHESIZED_WIRE_1610;
wire	SYNTHESIZED_WIRE_1611;
wire	SYNTHESIZED_WIRE_1612;
wire	SYNTHESIZED_WIRE_1613;
wire	SYNTHESIZED_WIRE_1614;
wire	SYNTHESIZED_WIRE_1615;
wire	SYNTHESIZED_WIRE_1616;
wire	SYNTHESIZED_WIRE_1617;
wire	SYNTHESIZED_WIRE_1618;
wire	SYNTHESIZED_WIRE_1619;
wire	SYNTHESIZED_WIRE_1620;
wire	SYNTHESIZED_WIRE_1621;
wire	SYNTHESIZED_WIRE_1622;
wire	SYNTHESIZED_WIRE_1623;
wire	SYNTHESIZED_WIRE_1624;
wire	SYNTHESIZED_WIRE_1625;
wire	SYNTHESIZED_WIRE_1626;
wire	SYNTHESIZED_WIRE_1627;
wire	SYNTHESIZED_WIRE_1628;
wire	SYNTHESIZED_WIRE_1629;
wire	SYNTHESIZED_WIRE_1630;
wire	SYNTHESIZED_WIRE_1631;
wire	SYNTHESIZED_WIRE_1632;
wire	SYNTHESIZED_WIRE_1633;
wire	SYNTHESIZED_WIRE_1634;
wire	SYNTHESIZED_WIRE_1635;
wire	SYNTHESIZED_WIRE_1636;
wire	SYNTHESIZED_WIRE_1637;
wire	SYNTHESIZED_WIRE_1638;
wire	SYNTHESIZED_WIRE_1639;
wire	SYNTHESIZED_WIRE_1640;
wire	SYNTHESIZED_WIRE_1641;
wire	SYNTHESIZED_WIRE_1642;
wire	SYNTHESIZED_WIRE_1643;
wire	SYNTHESIZED_WIRE_1644;
wire	SYNTHESIZED_WIRE_1645;
wire	SYNTHESIZED_WIRE_1646;
wire	SYNTHESIZED_WIRE_1647;
wire	SYNTHESIZED_WIRE_1648;
wire	SYNTHESIZED_WIRE_1649;
wire	SYNTHESIZED_WIRE_1650;
wire	SYNTHESIZED_WIRE_1651;
wire	SYNTHESIZED_WIRE_1652;
wire	SYNTHESIZED_WIRE_1653;
wire	SYNTHESIZED_WIRE_1654;
wire	SYNTHESIZED_WIRE_1655;
wire	SYNTHESIZED_WIRE_1656;
wire	SYNTHESIZED_WIRE_1657;
wire	SYNTHESIZED_WIRE_1658;
wire	SYNTHESIZED_WIRE_1659;
wire	SYNTHESIZED_WIRE_1660;
wire	SYNTHESIZED_WIRE_1661;
wire	SYNTHESIZED_WIRE_1662;
wire	SYNTHESIZED_WIRE_1663;
wire	SYNTHESIZED_WIRE_1664;
wire	SYNTHESIZED_WIRE_1665;
wire	SYNTHESIZED_WIRE_1666;
wire	SYNTHESIZED_WIRE_1667;
wire	SYNTHESIZED_WIRE_1668;
wire	SYNTHESIZED_WIRE_1669;
wire	SYNTHESIZED_WIRE_1670;
wire	SYNTHESIZED_WIRE_1671;
wire	SYNTHESIZED_WIRE_1672;
wire	SYNTHESIZED_WIRE_1673;
wire	SYNTHESIZED_WIRE_1674;
wire	SYNTHESIZED_WIRE_1675;
wire	SYNTHESIZED_WIRE_1676;
wire	SYNTHESIZED_WIRE_1677;
wire	SYNTHESIZED_WIRE_1678;
wire	SYNTHESIZED_WIRE_1679;
wire	SYNTHESIZED_WIRE_1680;
wire	SYNTHESIZED_WIRE_1681;
wire	SYNTHESIZED_WIRE_1682;
wire	SYNTHESIZED_WIRE_1683;
wire	SYNTHESIZED_WIRE_1684;
wire	SYNTHESIZED_WIRE_1685;
wire	SYNTHESIZED_WIRE_1686;
wire	SYNTHESIZED_WIRE_1687;
wire	SYNTHESIZED_WIRE_1688;
wire	SYNTHESIZED_WIRE_1689;
wire	SYNTHESIZED_WIRE_1690;
wire	SYNTHESIZED_WIRE_1691;
wire	SYNTHESIZED_WIRE_1692;
wire	SYNTHESIZED_WIRE_1693;
wire	SYNTHESIZED_WIRE_1694;
wire	SYNTHESIZED_WIRE_1695;
wire	SYNTHESIZED_WIRE_1696;
wire	SYNTHESIZED_WIRE_1697;
wire	SYNTHESIZED_WIRE_1698;
wire	SYNTHESIZED_WIRE_1699;
wire	SYNTHESIZED_WIRE_1700;
wire	SYNTHESIZED_WIRE_1701;
wire	SYNTHESIZED_WIRE_1702;
wire	SYNTHESIZED_WIRE_1703;
wire	SYNTHESIZED_WIRE_1704;
wire	SYNTHESIZED_WIRE_1705;
wire	SYNTHESIZED_WIRE_1706;
wire	SYNTHESIZED_WIRE_1707;
wire	SYNTHESIZED_WIRE_1708;
wire	SYNTHESIZED_WIRE_1709;
wire	SYNTHESIZED_WIRE_1710;
wire	SYNTHESIZED_WIRE_1711;
wire	SYNTHESIZED_WIRE_1712;
wire	SYNTHESIZED_WIRE_1713;
wire	SYNTHESIZED_WIRE_1714;
wire	SYNTHESIZED_WIRE_1715;
wire	SYNTHESIZED_WIRE_1716;
wire	SYNTHESIZED_WIRE_1717;
wire	SYNTHESIZED_WIRE_1718;
wire	SYNTHESIZED_WIRE_1719;
wire	SYNTHESIZED_WIRE_1720;
wire	SYNTHESIZED_WIRE_1721;
wire	SYNTHESIZED_WIRE_1722;
wire	SYNTHESIZED_WIRE_1723;
wire	SYNTHESIZED_WIRE_1724;
wire	SYNTHESIZED_WIRE_1725;
wire	SYNTHESIZED_WIRE_1726;
wire	SYNTHESIZED_WIRE_1727;
wire	SYNTHESIZED_WIRE_1728;
wire	SYNTHESIZED_WIRE_1729;
wire	SYNTHESIZED_WIRE_1730;
wire	SYNTHESIZED_WIRE_1731;
wire	SYNTHESIZED_WIRE_1732;
wire	SYNTHESIZED_WIRE_1733;
wire	SYNTHESIZED_WIRE_1734;
wire	SYNTHESIZED_WIRE_1735;
wire	SYNTHESIZED_WIRE_1736;
wire	SYNTHESIZED_WIRE_1737;
wire	SYNTHESIZED_WIRE_1738;
wire	SYNTHESIZED_WIRE_1739;
wire	SYNTHESIZED_WIRE_1740;
wire	SYNTHESIZED_WIRE_1741;
wire	SYNTHESIZED_WIRE_1742;
wire	SYNTHESIZED_WIRE_1743;
wire	SYNTHESIZED_WIRE_1744;
wire	SYNTHESIZED_WIRE_1745;
wire	SYNTHESIZED_WIRE_1746;
wire	SYNTHESIZED_WIRE_1747;
wire	SYNTHESIZED_WIRE_1748;
wire	SYNTHESIZED_WIRE_1749;
wire	SYNTHESIZED_WIRE_1750;
wire	SYNTHESIZED_WIRE_1751;
wire	SYNTHESIZED_WIRE_1752;
wire	SYNTHESIZED_WIRE_1753;
wire	SYNTHESIZED_WIRE_1754;
wire	SYNTHESIZED_WIRE_1755;
wire	SYNTHESIZED_WIRE_1756;
wire	SYNTHESIZED_WIRE_1757;
wire	SYNTHESIZED_WIRE_1758;
wire	SYNTHESIZED_WIRE_1759;
wire	SYNTHESIZED_WIRE_1760;
wire	SYNTHESIZED_WIRE_1761;
wire	SYNTHESIZED_WIRE_1762;
wire	SYNTHESIZED_WIRE_1763;
wire	SYNTHESIZED_WIRE_1764;
wire	SYNTHESIZED_WIRE_1765;
wire	SYNTHESIZED_WIRE_1766;
wire	SYNTHESIZED_WIRE_1767;
wire	SYNTHESIZED_WIRE_1768;
wire	SYNTHESIZED_WIRE_1769;
wire	SYNTHESIZED_WIRE_1770;
wire	SYNTHESIZED_WIRE_1771;
wire	SYNTHESIZED_WIRE_1772;
wire	SYNTHESIZED_WIRE_1773;
wire	SYNTHESIZED_WIRE_1774;
wire	SYNTHESIZED_WIRE_1775;
wire	SYNTHESIZED_WIRE_1776;
wire	SYNTHESIZED_WIRE_1777;
wire	SYNTHESIZED_WIRE_1778;
wire	SYNTHESIZED_WIRE_1779;
wire	SYNTHESIZED_WIRE_1780;
wire	SYNTHESIZED_WIRE_1781;
wire	SYNTHESIZED_WIRE_1782;
wire	SYNTHESIZED_WIRE_1783;
wire	SYNTHESIZED_WIRE_1784;
wire	SYNTHESIZED_WIRE_1785;
wire	SYNTHESIZED_WIRE_1786;
wire	SYNTHESIZED_WIRE_1787;
wire	SYNTHESIZED_WIRE_1788;
wire	SYNTHESIZED_WIRE_1789;
wire	SYNTHESIZED_WIRE_1790;
wire	SYNTHESIZED_WIRE_1791;
wire	SYNTHESIZED_WIRE_1792;
wire	SYNTHESIZED_WIRE_1793;
wire	SYNTHESIZED_WIRE_1794;
wire	SYNTHESIZED_WIRE_1795;
wire	SYNTHESIZED_WIRE_1796;
wire	SYNTHESIZED_WIRE_1797;
wire	SYNTHESIZED_WIRE_1798;
wire	SYNTHESIZED_WIRE_1799;
wire	SYNTHESIZED_WIRE_1800;
wire	SYNTHESIZED_WIRE_1801;
wire	SYNTHESIZED_WIRE_1802;
wire	SYNTHESIZED_WIRE_1803;
wire	SYNTHESIZED_WIRE_1804;
wire	SYNTHESIZED_WIRE_1805;
wire	SYNTHESIZED_WIRE_1806;
wire	SYNTHESIZED_WIRE_1807;
wire	SYNTHESIZED_WIRE_1808;
wire	SYNTHESIZED_WIRE_1809;
wire	SYNTHESIZED_WIRE_1810;
wire	SYNTHESIZED_WIRE_1811;
wire	SYNTHESIZED_WIRE_1812;
wire	SYNTHESIZED_WIRE_1813;
wire	SYNTHESIZED_WIRE_1814;
wire	SYNTHESIZED_WIRE_1815;
wire	SYNTHESIZED_WIRE_1816;
wire	SYNTHESIZED_WIRE_1817;
wire	SYNTHESIZED_WIRE_1818;
wire	SYNTHESIZED_WIRE_1819;
wire	SYNTHESIZED_WIRE_1820;
wire	SYNTHESIZED_WIRE_1821;
wire	SYNTHESIZED_WIRE_1822;
wire	SYNTHESIZED_WIRE_1823;
wire	SYNTHESIZED_WIRE_1824;
wire	SYNTHESIZED_WIRE_1825;
wire	SYNTHESIZED_WIRE_1826;
wire	SYNTHESIZED_WIRE_1827;
wire	SYNTHESIZED_WIRE_1828;
wire	SYNTHESIZED_WIRE_1829;
wire	SYNTHESIZED_WIRE_1830;
wire	SYNTHESIZED_WIRE_1831;
wire	SYNTHESIZED_WIRE_1832;
wire	SYNTHESIZED_WIRE_1833;
wire	SYNTHESIZED_WIRE_1834;
wire	SYNTHESIZED_WIRE_1835;
wire	SYNTHESIZED_WIRE_1836;
wire	SYNTHESIZED_WIRE_1837;
wire	SYNTHESIZED_WIRE_1838;
wire	SYNTHESIZED_WIRE_1839;
wire	SYNTHESIZED_WIRE_1840;
wire	SYNTHESIZED_WIRE_1841;
wire	SYNTHESIZED_WIRE_1842;
wire	SYNTHESIZED_WIRE_1843;
wire	SYNTHESIZED_WIRE_1844;
wire	SYNTHESIZED_WIRE_1845;
wire	SYNTHESIZED_WIRE_1846;
wire	SYNTHESIZED_WIRE_1847;
wire	SYNTHESIZED_WIRE_1848;
wire	SYNTHESIZED_WIRE_1849;
wire	SYNTHESIZED_WIRE_1850;
wire	SYNTHESIZED_WIRE_1851;
wire	SYNTHESIZED_WIRE_1852;
wire	SYNTHESIZED_WIRE_1853;
wire	SYNTHESIZED_WIRE_1854;
wire	SYNTHESIZED_WIRE_1855;
wire	SYNTHESIZED_WIRE_1856;
wire	SYNTHESIZED_WIRE_1857;
wire	SYNTHESIZED_WIRE_1858;
wire	SYNTHESIZED_WIRE_1859;
wire	SYNTHESIZED_WIRE_1860;
wire	SYNTHESIZED_WIRE_1861;
wire	SYNTHESIZED_WIRE_1862;
wire	SYNTHESIZED_WIRE_1863;
wire	SYNTHESIZED_WIRE_1864;
wire	SYNTHESIZED_WIRE_1865;
wire	SYNTHESIZED_WIRE_1866;
wire	SYNTHESIZED_WIRE_1867;
wire	SYNTHESIZED_WIRE_1868;
wire	SYNTHESIZED_WIRE_1869;
wire	SYNTHESIZED_WIRE_1870;
wire	SYNTHESIZED_WIRE_1871;
wire	SYNTHESIZED_WIRE_1872;
wire	SYNTHESIZED_WIRE_1873;
wire	SYNTHESIZED_WIRE_1874;
wire	SYNTHESIZED_WIRE_1875;
wire	SYNTHESIZED_WIRE_1876;
wire	SYNTHESIZED_WIRE_1877;
wire	SYNTHESIZED_WIRE_1878;
wire	SYNTHESIZED_WIRE_1879;
wire	SYNTHESIZED_WIRE_1880;
wire	SYNTHESIZED_WIRE_1881;
wire	SYNTHESIZED_WIRE_1882;
wire	SYNTHESIZED_WIRE_1883;
wire	SYNTHESIZED_WIRE_1884;
wire	SYNTHESIZED_WIRE_1885;
wire	SYNTHESIZED_WIRE_1886;
wire	SYNTHESIZED_WIRE_1887;
wire	SYNTHESIZED_WIRE_1888;
wire	SYNTHESIZED_WIRE_1889;
wire	SYNTHESIZED_WIRE_1890;
wire	SYNTHESIZED_WIRE_1891;
wire	SYNTHESIZED_WIRE_1892;
wire	SYNTHESIZED_WIRE_1893;
wire	SYNTHESIZED_WIRE_1894;
wire	SYNTHESIZED_WIRE_1895;
wire	SYNTHESIZED_WIRE_1896;
wire	SYNTHESIZED_WIRE_1897;
wire	SYNTHESIZED_WIRE_1898;
wire	SYNTHESIZED_WIRE_1899;
wire	SYNTHESIZED_WIRE_1900;
wire	SYNTHESIZED_WIRE_1901;
wire	SYNTHESIZED_WIRE_1902;
wire	SYNTHESIZED_WIRE_1903;
wire	SYNTHESIZED_WIRE_1904;
wire	SYNTHESIZED_WIRE_1905;
wire	SYNTHESIZED_WIRE_1906;
wire	SYNTHESIZED_WIRE_1907;
wire	SYNTHESIZED_WIRE_1908;
wire	SYNTHESIZED_WIRE_1909;
wire	SYNTHESIZED_WIRE_1910;
wire	SYNTHESIZED_WIRE_1911;
wire	SYNTHESIZED_WIRE_1912;
wire	SYNTHESIZED_WIRE_1913;
wire	SYNTHESIZED_WIRE_1914;
wire	SYNTHESIZED_WIRE_1915;
wire	SYNTHESIZED_WIRE_1916;
wire	SYNTHESIZED_WIRE_1917;
wire	SYNTHESIZED_WIRE_1918;
wire	SYNTHESIZED_WIRE_1919;
wire	SYNTHESIZED_WIRE_1920;
wire	SYNTHESIZED_WIRE_1921;
wire	SYNTHESIZED_WIRE_1922;
wire	SYNTHESIZED_WIRE_1923;
wire	SYNTHESIZED_WIRE_1924;
wire	SYNTHESIZED_WIRE_1925;
wire	SYNTHESIZED_WIRE_1926;
wire	SYNTHESIZED_WIRE_1927;
wire	SYNTHESIZED_WIRE_1928;
wire	SYNTHESIZED_WIRE_1929;
wire	SYNTHESIZED_WIRE_1930;
wire	SYNTHESIZED_WIRE_1931;
wire	SYNTHESIZED_WIRE_1932;
wire	SYNTHESIZED_WIRE_1933;
wire	SYNTHESIZED_WIRE_1934;
wire	SYNTHESIZED_WIRE_1935;
wire	SYNTHESIZED_WIRE_1936;
wire	SYNTHESIZED_WIRE_1937;
wire	SYNTHESIZED_WIRE_1938;
wire	SYNTHESIZED_WIRE_1939;
wire	SYNTHESIZED_WIRE_1940;
wire	SYNTHESIZED_WIRE_1941;
wire	SYNTHESIZED_WIRE_1942;
wire	SYNTHESIZED_WIRE_1943;
wire	SYNTHESIZED_WIRE_1944;
wire	SYNTHESIZED_WIRE_1945;
wire	SYNTHESIZED_WIRE_1946;
wire	SYNTHESIZED_WIRE_1947;
wire	SYNTHESIZED_WIRE_1948;
wire	SYNTHESIZED_WIRE_1949;
wire	SYNTHESIZED_WIRE_1950;
wire	SYNTHESIZED_WIRE_1951;
wire	SYNTHESIZED_WIRE_1952;
wire	SYNTHESIZED_WIRE_1953;
wire	SYNTHESIZED_WIRE_1954;
wire	SYNTHESIZED_WIRE_1955;
wire	SYNTHESIZED_WIRE_1956;
wire	SYNTHESIZED_WIRE_1957;
wire	SYNTHESIZED_WIRE_1958;
wire	SYNTHESIZED_WIRE_1959;
wire	SYNTHESIZED_WIRE_1960;
wire	SYNTHESIZED_WIRE_1961;
wire	SYNTHESIZED_WIRE_1962;
wire	SYNTHESIZED_WIRE_1963;
wire	SYNTHESIZED_WIRE_1964;
wire	SYNTHESIZED_WIRE_1965;
wire	SYNTHESIZED_WIRE_1966;
wire	SYNTHESIZED_WIRE_1967;
wire	SYNTHESIZED_WIRE_1968;
wire	SYNTHESIZED_WIRE_1969;
wire	SYNTHESIZED_WIRE_1970;
wire	SYNTHESIZED_WIRE_1971;
wire	SYNTHESIZED_WIRE_1972;
wire	SYNTHESIZED_WIRE_1973;
wire	SYNTHESIZED_WIRE_1974;
wire	SYNTHESIZED_WIRE_1975;
wire	SYNTHESIZED_WIRE_1976;
wire	SYNTHESIZED_WIRE_1977;
wire	SYNTHESIZED_WIRE_1978;
wire	SYNTHESIZED_WIRE_1979;
wire	SYNTHESIZED_WIRE_1980;
wire	SYNTHESIZED_WIRE_1981;
wire	SYNTHESIZED_WIRE_1982;
wire	SYNTHESIZED_WIRE_1983;
wire	SYNTHESIZED_WIRE_1984;
wire	SYNTHESIZED_WIRE_1985;
wire	SYNTHESIZED_WIRE_1986;
wire	SYNTHESIZED_WIRE_1987;
wire	SYNTHESIZED_WIRE_1988;
wire	SYNTHESIZED_WIRE_1989;
wire	SYNTHESIZED_WIRE_1990;
wire	SYNTHESIZED_WIRE_1991;
wire	SYNTHESIZED_WIRE_1992;
wire	SYNTHESIZED_WIRE_1993;
wire	SYNTHESIZED_WIRE_1994;
wire	SYNTHESIZED_WIRE_1995;
wire	SYNTHESIZED_WIRE_1996;
wire	SYNTHESIZED_WIRE_1997;
wire	SYNTHESIZED_WIRE_1998;
wire	SYNTHESIZED_WIRE_1999;
wire	SYNTHESIZED_WIRE_2000;
wire	SYNTHESIZED_WIRE_2001;
wire	SYNTHESIZED_WIRE_2002;
wire	SYNTHESIZED_WIRE_2003;
wire	SYNTHESIZED_WIRE_2004;
wire	SYNTHESIZED_WIRE_2005;
wire	SYNTHESIZED_WIRE_2006;
wire	SYNTHESIZED_WIRE_2007;
wire	SYNTHESIZED_WIRE_2008;
wire	SYNTHESIZED_WIRE_2009;
wire	SYNTHESIZED_WIRE_2010;
wire	SYNTHESIZED_WIRE_2011;
wire	SYNTHESIZED_WIRE_2012;
wire	SYNTHESIZED_WIRE_2013;
wire	SYNTHESIZED_WIRE_2014;
wire	SYNTHESIZED_WIRE_2015;
wire	SYNTHESIZED_WIRE_2016;
wire	SYNTHESIZED_WIRE_2017;
wire	SYNTHESIZED_WIRE_2018;
wire	SYNTHESIZED_WIRE_2019;
wire	SYNTHESIZED_WIRE_2020;
wire	SYNTHESIZED_WIRE_2021;
wire	SYNTHESIZED_WIRE_2022;
wire	SYNTHESIZED_WIRE_2023;
wire	SYNTHESIZED_WIRE_2024;
wire	SYNTHESIZED_WIRE_2025;
wire	SYNTHESIZED_WIRE_2026;
wire	SYNTHESIZED_WIRE_2027;
wire	SYNTHESIZED_WIRE_2028;
wire	SYNTHESIZED_WIRE_2029;
wire	SYNTHESIZED_WIRE_2030;
wire	SYNTHESIZED_WIRE_2031;
wire	SYNTHESIZED_WIRE_2032;
wire	SYNTHESIZED_WIRE_2033;
wire	SYNTHESIZED_WIRE_2034;
wire	SYNTHESIZED_WIRE_2035;
wire	SYNTHESIZED_WIRE_2036;
wire	SYNTHESIZED_WIRE_2037;
wire	SYNTHESIZED_WIRE_2038;
wire	SYNTHESIZED_WIRE_2039;
wire	SYNTHESIZED_WIRE_2040;
wire	SYNTHESIZED_WIRE_2041;
wire	SYNTHESIZED_WIRE_2042;
wire	SYNTHESIZED_WIRE_2043;
wire	SYNTHESIZED_WIRE_2044;
wire	SYNTHESIZED_WIRE_2045;
wire	SYNTHESIZED_WIRE_2046;
wire	SYNTHESIZED_WIRE_2047;
wire	SYNTHESIZED_WIRE_2048;
wire	SYNTHESIZED_WIRE_2049;
wire	SYNTHESIZED_WIRE_2050;
wire	SYNTHESIZED_WIRE_2051;
wire	SYNTHESIZED_WIRE_2052;
wire	SYNTHESIZED_WIRE_2053;
wire	SYNTHESIZED_WIRE_2054;
wire	SYNTHESIZED_WIRE_2055;
wire	SYNTHESIZED_WIRE_2056;
wire	SYNTHESIZED_WIRE_2057;
wire	SYNTHESIZED_WIRE_2058;
wire	SYNTHESIZED_WIRE_2059;
wire	SYNTHESIZED_WIRE_2060;
wire	SYNTHESIZED_WIRE_2061;
wire	SYNTHESIZED_WIRE_2062;
wire	SYNTHESIZED_WIRE_2063;
wire	SYNTHESIZED_WIRE_2064;
wire	SYNTHESIZED_WIRE_2065;
wire	SYNTHESIZED_WIRE_2066;
wire	SYNTHESIZED_WIRE_2067;
wire	SYNTHESIZED_WIRE_2068;
wire	SYNTHESIZED_WIRE_2069;
wire	SYNTHESIZED_WIRE_2070;
wire	SYNTHESIZED_WIRE_2071;
wire	SYNTHESIZED_WIRE_2072;
wire	SYNTHESIZED_WIRE_2073;
wire	SYNTHESIZED_WIRE_2074;
wire	SYNTHESIZED_WIRE_2075;
wire	SYNTHESIZED_WIRE_2076;
wire	SYNTHESIZED_WIRE_2077;
wire	SYNTHESIZED_WIRE_2078;
wire	SYNTHESIZED_WIRE_2079;
wire	SYNTHESIZED_WIRE_2080;
wire	SYNTHESIZED_WIRE_2081;
wire	SYNTHESIZED_WIRE_2082;
wire	SYNTHESIZED_WIRE_2083;
wire	SYNTHESIZED_WIRE_2084;
wire	SYNTHESIZED_WIRE_2085;
wire	SYNTHESIZED_WIRE_2086;
wire	SYNTHESIZED_WIRE_2087;
wire	SYNTHESIZED_WIRE_2088;
wire	SYNTHESIZED_WIRE_2089;
wire	SYNTHESIZED_WIRE_2090;
wire	SYNTHESIZED_WIRE_2091;
wire	SYNTHESIZED_WIRE_2092;
wire	SYNTHESIZED_WIRE_2093;
wire	SYNTHESIZED_WIRE_2094;
wire	SYNTHESIZED_WIRE_2095;
wire	SYNTHESIZED_WIRE_2096;
wire	SYNTHESIZED_WIRE_2097;
wire	SYNTHESIZED_WIRE_2098;
wire	SYNTHESIZED_WIRE_2099;
wire	SYNTHESIZED_WIRE_2100;
wire	SYNTHESIZED_WIRE_2101;
wire	SYNTHESIZED_WIRE_2102;
wire	SYNTHESIZED_WIRE_2103;
wire	SYNTHESIZED_WIRE_2104;
wire	SYNTHESIZED_WIRE_2105;
wire	SYNTHESIZED_WIRE_2106;
wire	SYNTHESIZED_WIRE_2107;
wire	SYNTHESIZED_WIRE_2108;
wire	SYNTHESIZED_WIRE_2109;
wire	SYNTHESIZED_WIRE_2110;
wire	SYNTHESIZED_WIRE_2111;
wire	SYNTHESIZED_WIRE_2112;
wire	SYNTHESIZED_WIRE_2113;
wire	SYNTHESIZED_WIRE_2114;
wire	SYNTHESIZED_WIRE_2115;
wire	SYNTHESIZED_WIRE_2116;
wire	SYNTHESIZED_WIRE_2117;
wire	SYNTHESIZED_WIRE_2118;
wire	SYNTHESIZED_WIRE_2119;
wire	SYNTHESIZED_WIRE_2120;
wire	SYNTHESIZED_WIRE_2121;
wire	SYNTHESIZED_WIRE_2122;
wire	SYNTHESIZED_WIRE_2123;
wire	SYNTHESIZED_WIRE_2124;
wire	SYNTHESIZED_WIRE_2125;
wire	SYNTHESIZED_WIRE_2126;
wire	SYNTHESIZED_WIRE_2127;
wire	SYNTHESIZED_WIRE_2128;
wire	SYNTHESIZED_WIRE_2129;
wire	SYNTHESIZED_WIRE_2130;
wire	SYNTHESIZED_WIRE_2131;
wire	SYNTHESIZED_WIRE_2132;
wire	SYNTHESIZED_WIRE_2133;
wire	SYNTHESIZED_WIRE_2134;
wire	SYNTHESIZED_WIRE_2135;
wire	SYNTHESIZED_WIRE_2136;
wire	SYNTHESIZED_WIRE_2137;
wire	SYNTHESIZED_WIRE_2138;
wire	SYNTHESIZED_WIRE_2139;
wire	SYNTHESIZED_WIRE_2140;
wire	SYNTHESIZED_WIRE_2141;
wire	SYNTHESIZED_WIRE_2142;
wire	SYNTHESIZED_WIRE_2143;
wire	SYNTHESIZED_WIRE_2144;
wire	SYNTHESIZED_WIRE_2145;
wire	SYNTHESIZED_WIRE_2146;
wire	SYNTHESIZED_WIRE_2147;
wire	SYNTHESIZED_WIRE_2148;
wire	SYNTHESIZED_WIRE_2149;
wire	SYNTHESIZED_WIRE_2150;
wire	SYNTHESIZED_WIRE_2151;
wire	SYNTHESIZED_WIRE_2152;
wire	SYNTHESIZED_WIRE_2153;
wire	SYNTHESIZED_WIRE_2154;
wire	SYNTHESIZED_WIRE_2155;
wire	SYNTHESIZED_WIRE_2156;
wire	SYNTHESIZED_WIRE_2157;
wire	SYNTHESIZED_WIRE_2158;
wire	SYNTHESIZED_WIRE_2159;
wire	SYNTHESIZED_WIRE_2160;
wire	SYNTHESIZED_WIRE_2161;
wire	SYNTHESIZED_WIRE_2162;
wire	SYNTHESIZED_WIRE_2163;
wire	SYNTHESIZED_WIRE_2164;
wire	SYNTHESIZED_WIRE_2165;
wire	SYNTHESIZED_WIRE_2166;
wire	SYNTHESIZED_WIRE_2167;
wire	SYNTHESIZED_WIRE_2168;
wire	SYNTHESIZED_WIRE_2169;
wire	SYNTHESIZED_WIRE_2170;
wire	SYNTHESIZED_WIRE_2171;
wire	SYNTHESIZED_WIRE_2172;
wire	SYNTHESIZED_WIRE_2173;
wire	SYNTHESIZED_WIRE_2174;
wire	SYNTHESIZED_WIRE_2175;
wire	SYNTHESIZED_WIRE_2176;
wire	SYNTHESIZED_WIRE_2177;
wire	SYNTHESIZED_WIRE_2178;
wire	SYNTHESIZED_WIRE_2179;
wire	SYNTHESIZED_WIRE_2180;
wire	SYNTHESIZED_WIRE_2181;
wire	SYNTHESIZED_WIRE_2182;
wire	SYNTHESIZED_WIRE_2183;
wire	SYNTHESIZED_WIRE_2184;
wire	SYNTHESIZED_WIRE_2185;
wire	SYNTHESIZED_WIRE_2186;
wire	SYNTHESIZED_WIRE_2187;
wire	SYNTHESIZED_WIRE_2188;
wire	SYNTHESIZED_WIRE_2189;
wire	SYNTHESIZED_WIRE_2190;
wire	SYNTHESIZED_WIRE_2191;
wire	SYNTHESIZED_WIRE_2192;
wire	SYNTHESIZED_WIRE_2193;
wire	SYNTHESIZED_WIRE_2194;
wire	SYNTHESIZED_WIRE_2195;
wire	SYNTHESIZED_WIRE_2196;
wire	SYNTHESIZED_WIRE_2197;
wire	SYNTHESIZED_WIRE_2198;
wire	SYNTHESIZED_WIRE_2199;
wire	SYNTHESIZED_WIRE_2200;
wire	SYNTHESIZED_WIRE_2201;
wire	SYNTHESIZED_WIRE_2202;
wire	SYNTHESIZED_WIRE_2203;
wire	SYNTHESIZED_WIRE_2204;
wire	SYNTHESIZED_WIRE_2205;
wire	SYNTHESIZED_WIRE_2206;
wire	SYNTHESIZED_WIRE_2207;
wire	SYNTHESIZED_WIRE_2208;
wire	SYNTHESIZED_WIRE_2209;
wire	SYNTHESIZED_WIRE_2210;
wire	SYNTHESIZED_WIRE_2211;
wire	SYNTHESIZED_WIRE_2212;
wire	SYNTHESIZED_WIRE_2213;
wire	SYNTHESIZED_WIRE_2214;
wire	SYNTHESIZED_WIRE_2215;
wire	SYNTHESIZED_WIRE_2216;
wire	SYNTHESIZED_WIRE_2217;
wire	SYNTHESIZED_WIRE_2218;
wire	SYNTHESIZED_WIRE_2219;
wire	SYNTHESIZED_WIRE_2220;
wire	SYNTHESIZED_WIRE_2221;
wire	SYNTHESIZED_WIRE_2222;
wire	SYNTHESIZED_WIRE_2223;
wire	SYNTHESIZED_WIRE_2224;
wire	SYNTHESIZED_WIRE_2225;
wire	SYNTHESIZED_WIRE_2226;
wire	SYNTHESIZED_WIRE_2227;
wire	SYNTHESIZED_WIRE_2228;
wire	SYNTHESIZED_WIRE_2229;
wire	SYNTHESIZED_WIRE_2230;
wire	SYNTHESIZED_WIRE_2231;
wire	SYNTHESIZED_WIRE_2232;
wire	SYNTHESIZED_WIRE_2233;
wire	SYNTHESIZED_WIRE_2234;
wire	SYNTHESIZED_WIRE_2235;
wire	SYNTHESIZED_WIRE_2236;
wire	SYNTHESIZED_WIRE_2237;
wire	SYNTHESIZED_WIRE_2238;
wire	SYNTHESIZED_WIRE_2239;
wire	SYNTHESIZED_WIRE_2240;
wire	SYNTHESIZED_WIRE_2241;
wire	SYNTHESIZED_WIRE_2242;
wire	SYNTHESIZED_WIRE_2243;
wire	SYNTHESIZED_WIRE_2244;
wire	SYNTHESIZED_WIRE_2245;
wire	SYNTHESIZED_WIRE_2246;
wire	SYNTHESIZED_WIRE_2247;
wire	SYNTHESIZED_WIRE_2248;
wire	SYNTHESIZED_WIRE_2249;
wire	SYNTHESIZED_WIRE_2250;
wire	SYNTHESIZED_WIRE_2251;
wire	SYNTHESIZED_WIRE_2252;
wire	SYNTHESIZED_WIRE_2253;
wire	SYNTHESIZED_WIRE_2254;
wire	SYNTHESIZED_WIRE_2255;
wire	SYNTHESIZED_WIRE_2256;
wire	SYNTHESIZED_WIRE_2257;
wire	SYNTHESIZED_WIRE_2258;
wire	SYNTHESIZED_WIRE_2259;
wire	SYNTHESIZED_WIRE_2260;
wire	SYNTHESIZED_WIRE_2261;
wire	SYNTHESIZED_WIRE_2262;
wire	SYNTHESIZED_WIRE_2263;
wire	SYNTHESIZED_WIRE_2264;
wire	SYNTHESIZED_WIRE_2265;
wire	SYNTHESIZED_WIRE_2266;
wire	SYNTHESIZED_WIRE_2267;
wire	SYNTHESIZED_WIRE_2268;
wire	SYNTHESIZED_WIRE_2269;
wire	SYNTHESIZED_WIRE_2270;
wire	SYNTHESIZED_WIRE_2271;
wire	SYNTHESIZED_WIRE_2272;
wire	SYNTHESIZED_WIRE_2273;
wire	SYNTHESIZED_WIRE_2274;
wire	SYNTHESIZED_WIRE_2275;
wire	SYNTHESIZED_WIRE_2276;
wire	SYNTHESIZED_WIRE_2277;
wire	SYNTHESIZED_WIRE_2278;
wire	SYNTHESIZED_WIRE_2279;
wire	SYNTHESIZED_WIRE_2280;
wire	SYNTHESIZED_WIRE_2281;
wire	SYNTHESIZED_WIRE_2282;
wire	SYNTHESIZED_WIRE_2283;
wire	SYNTHESIZED_WIRE_2284;
wire	SYNTHESIZED_WIRE_2285;
wire	SYNTHESIZED_WIRE_2286;
wire	SYNTHESIZED_WIRE_2287;
wire	SYNTHESIZED_WIRE_2288;
wire	SYNTHESIZED_WIRE_2289;
wire	SYNTHESIZED_WIRE_2290;
wire	SYNTHESIZED_WIRE_2291;
wire	SYNTHESIZED_WIRE_2292;
wire	SYNTHESIZED_WIRE_2293;
wire	SYNTHESIZED_WIRE_2294;
wire	SYNTHESIZED_WIRE_2295;
wire	SYNTHESIZED_WIRE_2296;
wire	SYNTHESIZED_WIRE_2297;
wire	SYNTHESIZED_WIRE_2298;
wire	SYNTHESIZED_WIRE_2299;
wire	SYNTHESIZED_WIRE_2300;
wire	SYNTHESIZED_WIRE_2301;
wire	SYNTHESIZED_WIRE_2302;
wire	SYNTHESIZED_WIRE_2303;
wire	SYNTHESIZED_WIRE_2304;
wire	SYNTHESIZED_WIRE_2305;
wire	SYNTHESIZED_WIRE_2306;
wire	SYNTHESIZED_WIRE_2307;
wire	SYNTHESIZED_WIRE_2308;
wire	SYNTHESIZED_WIRE_2309;
wire	SYNTHESIZED_WIRE_2310;
wire	SYNTHESIZED_WIRE_2311;
wire	SYNTHESIZED_WIRE_2312;
wire	SYNTHESIZED_WIRE_2313;
wire	SYNTHESIZED_WIRE_2314;
wire	SYNTHESIZED_WIRE_2315;
wire	SYNTHESIZED_WIRE_2316;
wire	SYNTHESIZED_WIRE_2317;
wire	SYNTHESIZED_WIRE_2318;
wire	SYNTHESIZED_WIRE_2319;
wire	SYNTHESIZED_WIRE_2320;
wire	SYNTHESIZED_WIRE_2321;
wire	SYNTHESIZED_WIRE_2322;
wire	SYNTHESIZED_WIRE_2323;
wire	SYNTHESIZED_WIRE_2324;
wire	SYNTHESIZED_WIRE_2325;
wire	SYNTHESIZED_WIRE_2326;
wire	SYNTHESIZED_WIRE_2327;
wire	SYNTHESIZED_WIRE_2328;
wire	SYNTHESIZED_WIRE_2329;
wire	SYNTHESIZED_WIRE_2330;
wire	SYNTHESIZED_WIRE_2331;
wire	SYNTHESIZED_WIRE_2332;
wire	SYNTHESIZED_WIRE_2333;
wire	SYNTHESIZED_WIRE_2334;
wire	SYNTHESIZED_WIRE_2335;
wire	SYNTHESIZED_WIRE_2336;
wire	SYNTHESIZED_WIRE_2337;
wire	SYNTHESIZED_WIRE_2338;
wire	SYNTHESIZED_WIRE_2339;
wire	SYNTHESIZED_WIRE_2340;
wire	SYNTHESIZED_WIRE_2341;
wire	SYNTHESIZED_WIRE_2342;
wire	SYNTHESIZED_WIRE_2343;
wire	SYNTHESIZED_WIRE_2344;
wire	SYNTHESIZED_WIRE_2345;
wire	SYNTHESIZED_WIRE_2346;
wire	SYNTHESIZED_WIRE_2347;
wire	SYNTHESIZED_WIRE_2348;
wire	SYNTHESIZED_WIRE_2349;
wire	SYNTHESIZED_WIRE_2350;
wire	SYNTHESIZED_WIRE_2351;
wire	SYNTHESIZED_WIRE_2352;
wire	SYNTHESIZED_WIRE_2353;
wire	SYNTHESIZED_WIRE_2354;
wire	SYNTHESIZED_WIRE_2355;
wire	SYNTHESIZED_WIRE_2356;
wire	SYNTHESIZED_WIRE_2357;
wire	SYNTHESIZED_WIRE_2358;
wire	SYNTHESIZED_WIRE_2359;
wire	SYNTHESIZED_WIRE_2360;
wire	SYNTHESIZED_WIRE_2361;
wire	SYNTHESIZED_WIRE_2362;
wire	SYNTHESIZED_WIRE_2363;
wire	SYNTHESIZED_WIRE_2364;
wire	SYNTHESIZED_WIRE_2365;
wire	SYNTHESIZED_WIRE_2366;
wire	SYNTHESIZED_WIRE_2367;
wire	SYNTHESIZED_WIRE_2368;
wire	SYNTHESIZED_WIRE_2369;
wire	SYNTHESIZED_WIRE_2370;
wire	SYNTHESIZED_WIRE_2371;
wire	SYNTHESIZED_WIRE_2372;
wire	SYNTHESIZED_WIRE_2373;
wire	SYNTHESIZED_WIRE_2374;
wire	SYNTHESIZED_WIRE_2375;
wire	SYNTHESIZED_WIRE_2376;
wire	SYNTHESIZED_WIRE_2377;
wire	SYNTHESIZED_WIRE_2378;
wire	SYNTHESIZED_WIRE_2379;
wire	SYNTHESIZED_WIRE_2380;
wire	SYNTHESIZED_WIRE_2381;
wire	SYNTHESIZED_WIRE_2382;
wire	SYNTHESIZED_WIRE_2383;
wire	SYNTHESIZED_WIRE_2384;
wire	SYNTHESIZED_WIRE_2385;
wire	SYNTHESIZED_WIRE_2386;
wire	SYNTHESIZED_WIRE_2387;
wire	SYNTHESIZED_WIRE_2388;
wire	SYNTHESIZED_WIRE_2389;
wire	SYNTHESIZED_WIRE_2390;
wire	SYNTHESIZED_WIRE_2391;
wire	SYNTHESIZED_WIRE_2392;
wire	SYNTHESIZED_WIRE_2393;
wire	SYNTHESIZED_WIRE_2394;
wire	SYNTHESIZED_WIRE_2395;
wire	SYNTHESIZED_WIRE_2396;
wire	SYNTHESIZED_WIRE_2397;
wire	SYNTHESIZED_WIRE_2398;
wire	SYNTHESIZED_WIRE_2399;
wire	SYNTHESIZED_WIRE_2400;
wire	SYNTHESIZED_WIRE_2401;
wire	SYNTHESIZED_WIRE_2402;
wire	SYNTHESIZED_WIRE_2403;
wire	SYNTHESIZED_WIRE_2404;
wire	SYNTHESIZED_WIRE_2405;
wire	SYNTHESIZED_WIRE_2406;
wire	SYNTHESIZED_WIRE_2407;
wire	SYNTHESIZED_WIRE_2408;
wire	SYNTHESIZED_WIRE_2409;
wire	SYNTHESIZED_WIRE_2410;
wire	SYNTHESIZED_WIRE_2411;
wire	SYNTHESIZED_WIRE_2412;
wire	SYNTHESIZED_WIRE_2413;
wire	SYNTHESIZED_WIRE_2414;
wire	SYNTHESIZED_WIRE_2415;
wire	SYNTHESIZED_WIRE_2416;
wire	SYNTHESIZED_WIRE_2417;
wire	SYNTHESIZED_WIRE_2418;
wire	SYNTHESIZED_WIRE_2419;
wire	SYNTHESIZED_WIRE_2420;
wire	SYNTHESIZED_WIRE_2421;
wire	SYNTHESIZED_WIRE_2422;
wire	SYNTHESIZED_WIRE_2423;
wire	SYNTHESIZED_WIRE_2424;
wire	SYNTHESIZED_WIRE_2425;
wire	SYNTHESIZED_WIRE_2426;
wire	SYNTHESIZED_WIRE_2427;
wire	SYNTHESIZED_WIRE_2428;
wire	SYNTHESIZED_WIRE_2429;
wire	SYNTHESIZED_WIRE_2430;
wire	SYNTHESIZED_WIRE_2431;
wire	SYNTHESIZED_WIRE_2432;
wire	SYNTHESIZED_WIRE_2433;
wire	SYNTHESIZED_WIRE_2434;
wire	SYNTHESIZED_WIRE_2435;
wire	SYNTHESIZED_WIRE_2436;
wire	SYNTHESIZED_WIRE_2437;
wire	SYNTHESIZED_WIRE_2438;
wire	SYNTHESIZED_WIRE_2439;
wire	SYNTHESIZED_WIRE_2440;
wire	SYNTHESIZED_WIRE_2441;
wire	SYNTHESIZED_WIRE_2442;
wire	SYNTHESIZED_WIRE_2443;
wire	SYNTHESIZED_WIRE_2444;
wire	SYNTHESIZED_WIRE_2445;
wire	SYNTHESIZED_WIRE_2446;
wire	SYNTHESIZED_WIRE_2447;
wire	SYNTHESIZED_WIRE_2448;
wire	SYNTHESIZED_WIRE_2449;
wire	SYNTHESIZED_WIRE_2450;
wire	SYNTHESIZED_WIRE_2451;
wire	SYNTHESIZED_WIRE_2452;
wire	SYNTHESIZED_WIRE_2453;
wire	SYNTHESIZED_WIRE_2454;
wire	SYNTHESIZED_WIRE_2455;
wire	SYNTHESIZED_WIRE_2456;
wire	SYNTHESIZED_WIRE_2457;
wire	SYNTHESIZED_WIRE_2458;
wire	SYNTHESIZED_WIRE_2459;
wire	SYNTHESIZED_WIRE_2460;
wire	SYNTHESIZED_WIRE_2461;
wire	SYNTHESIZED_WIRE_2462;
wire	SYNTHESIZED_WIRE_2463;
wire	SYNTHESIZED_WIRE_2464;
wire	SYNTHESIZED_WIRE_2465;
wire	SYNTHESIZED_WIRE_2466;
wire	SYNTHESIZED_WIRE_2467;
wire	SYNTHESIZED_WIRE_2468;
wire	SYNTHESIZED_WIRE_2469;
wire	SYNTHESIZED_WIRE_2470;
wire	SYNTHESIZED_WIRE_2471;
wire	SYNTHESIZED_WIRE_2472;
wire	SYNTHESIZED_WIRE_2473;
wire	SYNTHESIZED_WIRE_2474;
wire	SYNTHESIZED_WIRE_2475;
wire	SYNTHESIZED_WIRE_2476;
wire	SYNTHESIZED_WIRE_2477;
wire	SYNTHESIZED_WIRE_2478;
wire	SYNTHESIZED_WIRE_2479;
wire	SYNTHESIZED_WIRE_2480;
wire	SYNTHESIZED_WIRE_2481;
wire	SYNTHESIZED_WIRE_2482;
wire	SYNTHESIZED_WIRE_2483;
wire	SYNTHESIZED_WIRE_2484;
wire	SYNTHESIZED_WIRE_2485;
wire	SYNTHESIZED_WIRE_2486;
wire	SYNTHESIZED_WIRE_2487;
wire	SYNTHESIZED_WIRE_2488;
wire	SYNTHESIZED_WIRE_2489;
wire	SYNTHESIZED_WIRE_2490;
wire	SYNTHESIZED_WIRE_2491;
wire	SYNTHESIZED_WIRE_2492;
wire	SYNTHESIZED_WIRE_2493;
wire	SYNTHESIZED_WIRE_2494;
wire	SYNTHESIZED_WIRE_2495;
wire	SYNTHESIZED_WIRE_2496;
wire	SYNTHESIZED_WIRE_2497;
wire	SYNTHESIZED_WIRE_2498;
wire	SYNTHESIZED_WIRE_2499;
wire	SYNTHESIZED_WIRE_2500;
wire	SYNTHESIZED_WIRE_2501;
wire	SYNTHESIZED_WIRE_2502;
wire	SYNTHESIZED_WIRE_2503;
wire	SYNTHESIZED_WIRE_2504;
wire	SYNTHESIZED_WIRE_2505;
wire	SYNTHESIZED_WIRE_2506;
wire	SYNTHESIZED_WIRE_2507;
wire	SYNTHESIZED_WIRE_2508;
wire	SYNTHESIZED_WIRE_2509;
wire	SYNTHESIZED_WIRE_2510;
wire	SYNTHESIZED_WIRE_2511;
wire	SYNTHESIZED_WIRE_2512;
wire	SYNTHESIZED_WIRE_2513;
wire	SYNTHESIZED_WIRE_2514;
wire	SYNTHESIZED_WIRE_2515;
wire	SYNTHESIZED_WIRE_2516;
wire	SYNTHESIZED_WIRE_2517;
wire	SYNTHESIZED_WIRE_2518;
wire	SYNTHESIZED_WIRE_2519;
wire	SYNTHESIZED_WIRE_2520;
wire	SYNTHESIZED_WIRE_2521;
wire	SYNTHESIZED_WIRE_2522;
wire	SYNTHESIZED_WIRE_2523;
wire	SYNTHESIZED_WIRE_2524;
wire	SYNTHESIZED_WIRE_2525;
wire	SYNTHESIZED_WIRE_2526;
wire	SYNTHESIZED_WIRE_2527;
wire	SYNTHESIZED_WIRE_2528;
wire	SYNTHESIZED_WIRE_2529;
wire	SYNTHESIZED_WIRE_2530;
wire	SYNTHESIZED_WIRE_2531;
wire	SYNTHESIZED_WIRE_2532;
wire	SYNTHESIZED_WIRE_2533;
wire	SYNTHESIZED_WIRE_2534;
wire	SYNTHESIZED_WIRE_2535;
wire	SYNTHESIZED_WIRE_2536;
wire	SYNTHESIZED_WIRE_2537;
wire	SYNTHESIZED_WIRE_2538;
wire	SYNTHESIZED_WIRE_2539;
wire	SYNTHESIZED_WIRE_2540;
wire	SYNTHESIZED_WIRE_2541;
wire	SYNTHESIZED_WIRE_2542;
wire	SYNTHESIZED_WIRE_2543;
wire	SYNTHESIZED_WIRE_2544;
wire	SYNTHESIZED_WIRE_2545;
wire	SYNTHESIZED_WIRE_2546;
wire	SYNTHESIZED_WIRE_2547;
wire	SYNTHESIZED_WIRE_2548;
wire	SYNTHESIZED_WIRE_2549;
wire	SYNTHESIZED_WIRE_2550;
wire	SYNTHESIZED_WIRE_2551;
wire	SYNTHESIZED_WIRE_2552;
wire	SYNTHESIZED_WIRE_2553;
wire	SYNTHESIZED_WIRE_2554;
wire	SYNTHESIZED_WIRE_2555;
wire	SYNTHESIZED_WIRE_2556;
wire	SYNTHESIZED_WIRE_2557;
wire	SYNTHESIZED_WIRE_2558;
wire	SYNTHESIZED_WIRE_2559;
wire	SYNTHESIZED_WIRE_2560;
wire	SYNTHESIZED_WIRE_2561;
wire	SYNTHESIZED_WIRE_2562;
wire	SYNTHESIZED_WIRE_2563;
wire	SYNTHESIZED_WIRE_2564;
wire	SYNTHESIZED_WIRE_2565;
wire	SYNTHESIZED_WIRE_2566;
wire	SYNTHESIZED_WIRE_2567;
wire	SYNTHESIZED_WIRE_2568;
wire	SYNTHESIZED_WIRE_2569;
wire	SYNTHESIZED_WIRE_2570;
wire	SYNTHESIZED_WIRE_2571;
wire	SYNTHESIZED_WIRE_2572;
wire	SYNTHESIZED_WIRE_2573;
wire	SYNTHESIZED_WIRE_2574;
wire	SYNTHESIZED_WIRE_2575;
wire	SYNTHESIZED_WIRE_2576;
wire	SYNTHESIZED_WIRE_2577;
wire	SYNTHESIZED_WIRE_2578;
wire	SYNTHESIZED_WIRE_2579;
wire	SYNTHESIZED_WIRE_2580;
wire	SYNTHESIZED_WIRE_2581;
wire	SYNTHESIZED_WIRE_2582;
wire	SYNTHESIZED_WIRE_2583;
wire	SYNTHESIZED_WIRE_2584;
wire	SYNTHESIZED_WIRE_2585;
wire	SYNTHESIZED_WIRE_2586;
wire	SYNTHESIZED_WIRE_2587;
wire	SYNTHESIZED_WIRE_2588;
wire	SYNTHESIZED_WIRE_2589;
wire	SYNTHESIZED_WIRE_2590;
wire	SYNTHESIZED_WIRE_2591;
wire	SYNTHESIZED_WIRE_2592;
wire	SYNTHESIZED_WIRE_2593;
wire	SYNTHESIZED_WIRE_2594;
wire	SYNTHESIZED_WIRE_2595;
wire	SYNTHESIZED_WIRE_2596;
wire	SYNTHESIZED_WIRE_2597;
wire	SYNTHESIZED_WIRE_2598;
wire	SYNTHESIZED_WIRE_2599;
wire	SYNTHESIZED_WIRE_2600;
wire	SYNTHESIZED_WIRE_2601;
wire	SYNTHESIZED_WIRE_2602;
wire	SYNTHESIZED_WIRE_2603;
wire	SYNTHESIZED_WIRE_2604;
wire	SYNTHESIZED_WIRE_2605;
wire	SYNTHESIZED_WIRE_2606;
wire	SYNTHESIZED_WIRE_2607;
wire	SYNTHESIZED_WIRE_2608;
wire	SYNTHESIZED_WIRE_2609;
wire	SYNTHESIZED_WIRE_2610;
wire	SYNTHESIZED_WIRE_2611;
wire	SYNTHESIZED_WIRE_2612;
wire	SYNTHESIZED_WIRE_2613;
wire	SYNTHESIZED_WIRE_2614;
wire	SYNTHESIZED_WIRE_2615;
wire	SYNTHESIZED_WIRE_2616;
wire	SYNTHESIZED_WIRE_2617;
wire	SYNTHESIZED_WIRE_2618;
wire	SYNTHESIZED_WIRE_2619;
wire	SYNTHESIZED_WIRE_2620;
wire	SYNTHESIZED_WIRE_2621;
wire	SYNTHESIZED_WIRE_2622;
wire	SYNTHESIZED_WIRE_2623;
wire	SYNTHESIZED_WIRE_2624;
wire	SYNTHESIZED_WIRE_2625;
wire	SYNTHESIZED_WIRE_2626;
wire	SYNTHESIZED_WIRE_2627;
wire	SYNTHESIZED_WIRE_2628;
wire	SYNTHESIZED_WIRE_2629;
wire	SYNTHESIZED_WIRE_2630;
wire	SYNTHESIZED_WIRE_2631;
wire	SYNTHESIZED_WIRE_2632;
wire	SYNTHESIZED_WIRE_2633;
wire	SYNTHESIZED_WIRE_2634;
wire	SYNTHESIZED_WIRE_2635;
wire	SYNTHESIZED_WIRE_2636;
wire	SYNTHESIZED_WIRE_2637;
wire	SYNTHESIZED_WIRE_2638;
wire	SYNTHESIZED_WIRE_2639;
wire	SYNTHESIZED_WIRE_2640;
wire	SYNTHESIZED_WIRE_2641;
wire	SYNTHESIZED_WIRE_2642;
wire	SYNTHESIZED_WIRE_2643;
wire	SYNTHESIZED_WIRE_2644;
wire	SYNTHESIZED_WIRE_2645;
wire	SYNTHESIZED_WIRE_2646;
wire	SYNTHESIZED_WIRE_2647;
wire	SYNTHESIZED_WIRE_2648;
wire	SYNTHESIZED_WIRE_2649;
wire	SYNTHESIZED_WIRE_2650;
wire	SYNTHESIZED_WIRE_2651;
wire	SYNTHESIZED_WIRE_2652;
wire	SYNTHESIZED_WIRE_2653;
wire	SYNTHESIZED_WIRE_2654;
wire	SYNTHESIZED_WIRE_2655;
wire	SYNTHESIZED_WIRE_2656;
wire	SYNTHESIZED_WIRE_2657;
wire	SYNTHESIZED_WIRE_2658;
wire	SYNTHESIZED_WIRE_2659;
wire	SYNTHESIZED_WIRE_2660;
wire	SYNTHESIZED_WIRE_2661;
wire	SYNTHESIZED_WIRE_2662;
wire	SYNTHESIZED_WIRE_2663;
wire	SYNTHESIZED_WIRE_2664;
wire	SYNTHESIZED_WIRE_2665;
wire	SYNTHESIZED_WIRE_2666;
wire	SYNTHESIZED_WIRE_2667;
wire	SYNTHESIZED_WIRE_2668;
wire	SYNTHESIZED_WIRE_2669;
wire	SYNTHESIZED_WIRE_2670;
wire	SYNTHESIZED_WIRE_2671;
wire	SYNTHESIZED_WIRE_2672;
wire	SYNTHESIZED_WIRE_2673;
wire	SYNTHESIZED_WIRE_2674;
wire	SYNTHESIZED_WIRE_2675;
wire	SYNTHESIZED_WIRE_2676;
wire	SYNTHESIZED_WIRE_2677;
wire	SYNTHESIZED_WIRE_2678;
wire	SYNTHESIZED_WIRE_2679;
wire	SYNTHESIZED_WIRE_2680;
wire	SYNTHESIZED_WIRE_2681;
wire	SYNTHESIZED_WIRE_2682;
wire	SYNTHESIZED_WIRE_2683;
wire	SYNTHESIZED_WIRE_2684;
wire	SYNTHESIZED_WIRE_2685;
wire	SYNTHESIZED_WIRE_2686;
wire	SYNTHESIZED_WIRE_2687;
wire	SYNTHESIZED_WIRE_2688;
wire	SYNTHESIZED_WIRE_2689;
wire	SYNTHESIZED_WIRE_2690;
wire	SYNTHESIZED_WIRE_2691;
wire	SYNTHESIZED_WIRE_2692;
wire	SYNTHESIZED_WIRE_2693;
wire	SYNTHESIZED_WIRE_2694;
wire	SYNTHESIZED_WIRE_2695;
wire	SYNTHESIZED_WIRE_2696;
wire	SYNTHESIZED_WIRE_2697;
wire	SYNTHESIZED_WIRE_2698;
wire	SYNTHESIZED_WIRE_2699;
wire	SYNTHESIZED_WIRE_2700;
wire	SYNTHESIZED_WIRE_2701;
wire	SYNTHESIZED_WIRE_2702;
wire	SYNTHESIZED_WIRE_2703;
wire	SYNTHESIZED_WIRE_2704;
wire	SYNTHESIZED_WIRE_2705;
wire	SYNTHESIZED_WIRE_2706;
wire	SYNTHESIZED_WIRE_2707;
wire	SYNTHESIZED_WIRE_2708;
wire	SYNTHESIZED_WIRE_2709;
wire	SYNTHESIZED_WIRE_2710;
wire	SYNTHESIZED_WIRE_2711;
wire	SYNTHESIZED_WIRE_2712;
wire	SYNTHESIZED_WIRE_2713;
wire	SYNTHESIZED_WIRE_2714;
wire	SYNTHESIZED_WIRE_2715;
wire	SYNTHESIZED_WIRE_2716;
wire	SYNTHESIZED_WIRE_2717;
wire	SYNTHESIZED_WIRE_2718;
wire	SYNTHESIZED_WIRE_2719;
wire	SYNTHESIZED_WIRE_2720;
wire	SYNTHESIZED_WIRE_2721;
wire	SYNTHESIZED_WIRE_2722;
wire	SYNTHESIZED_WIRE_2723;
wire	SYNTHESIZED_WIRE_2724;
wire	SYNTHESIZED_WIRE_2725;
wire	SYNTHESIZED_WIRE_2726;
wire	SYNTHESIZED_WIRE_2727;
wire	SYNTHESIZED_WIRE_2728;
wire	SYNTHESIZED_WIRE_2729;
wire	SYNTHESIZED_WIRE_2730;
wire	SYNTHESIZED_WIRE_2731;
wire	SYNTHESIZED_WIRE_2732;
wire	SYNTHESIZED_WIRE_2733;
wire	SYNTHESIZED_WIRE_2734;
wire	SYNTHESIZED_WIRE_2735;
wire	SYNTHESIZED_WIRE_2736;
wire	SYNTHESIZED_WIRE_2737;
wire	SYNTHESIZED_WIRE_2738;
wire	SYNTHESIZED_WIRE_2739;
wire	SYNTHESIZED_WIRE_2740;
wire	SYNTHESIZED_WIRE_2741;
wire	SYNTHESIZED_WIRE_2742;
wire	SYNTHESIZED_WIRE_2743;
wire	SYNTHESIZED_WIRE_2744;
wire	SYNTHESIZED_WIRE_2745;
wire	SYNTHESIZED_WIRE_2746;
wire	SYNTHESIZED_WIRE_2747;
wire	SYNTHESIZED_WIRE_2748;
wire	SYNTHESIZED_WIRE_2749;
wire	SYNTHESIZED_WIRE_2750;
wire	SYNTHESIZED_WIRE_2751;
wire	SYNTHESIZED_WIRE_2752;
wire	SYNTHESIZED_WIRE_2753;
wire	SYNTHESIZED_WIRE_2754;
wire	SYNTHESIZED_WIRE_2755;
wire	SYNTHESIZED_WIRE_2756;
wire	SYNTHESIZED_WIRE_2757;
wire	SYNTHESIZED_WIRE_2758;
wire	SYNTHESIZED_WIRE_2759;
wire	SYNTHESIZED_WIRE_2760;
wire	SYNTHESIZED_WIRE_2761;
wire	SYNTHESIZED_WIRE_2762;
wire	SYNTHESIZED_WIRE_2763;
wire	SYNTHESIZED_WIRE_2764;
wire	SYNTHESIZED_WIRE_2765;
wire	SYNTHESIZED_WIRE_2766;
wire	SYNTHESIZED_WIRE_2767;
wire	SYNTHESIZED_WIRE_2768;
wire	SYNTHESIZED_WIRE_2769;
wire	SYNTHESIZED_WIRE_2770;
wire	SYNTHESIZED_WIRE_2771;
wire	SYNTHESIZED_WIRE_2772;
wire	SYNTHESIZED_WIRE_2773;
wire	SYNTHESIZED_WIRE_2774;
wire	SYNTHESIZED_WIRE_2775;
wire	SYNTHESIZED_WIRE_2776;
wire	SYNTHESIZED_WIRE_2777;
wire	SYNTHESIZED_WIRE_2778;
wire	SYNTHESIZED_WIRE_2779;
wire	SYNTHESIZED_WIRE_2780;
wire	SYNTHESIZED_WIRE_2781;
wire	SYNTHESIZED_WIRE_2782;
wire	SYNTHESIZED_WIRE_2783;
wire	SYNTHESIZED_WIRE_2784;
wire	SYNTHESIZED_WIRE_2785;
wire	SYNTHESIZED_WIRE_2786;
wire	SYNTHESIZED_WIRE_2787;
wire	SYNTHESIZED_WIRE_2788;
wire	SYNTHESIZED_WIRE_2789;
wire	SYNTHESIZED_WIRE_2790;
wire	SYNTHESIZED_WIRE_2791;
wire	SYNTHESIZED_WIRE_2792;
wire	SYNTHESIZED_WIRE_2793;
wire	SYNTHESIZED_WIRE_2794;
wire	SYNTHESIZED_WIRE_2795;
wire	SYNTHESIZED_WIRE_2796;
wire	SYNTHESIZED_WIRE_2797;
wire	SYNTHESIZED_WIRE_2798;
wire	SYNTHESIZED_WIRE_2799;
wire	SYNTHESIZED_WIRE_2800;
wire	SYNTHESIZED_WIRE_2801;
wire	SYNTHESIZED_WIRE_2802;
wire	SYNTHESIZED_WIRE_2803;
wire	SYNTHESIZED_WIRE_2804;
wire	SYNTHESIZED_WIRE_2805;
wire	SYNTHESIZED_WIRE_2806;
wire	SYNTHESIZED_WIRE_2807;
wire	SYNTHESIZED_WIRE_2808;
wire	SYNTHESIZED_WIRE_2809;
wire	SYNTHESIZED_WIRE_2810;
wire	SYNTHESIZED_WIRE_2811;
wire	SYNTHESIZED_WIRE_2812;
wire	SYNTHESIZED_WIRE_2813;
wire	SYNTHESIZED_WIRE_2814;
wire	SYNTHESIZED_WIRE_2815;
wire	SYNTHESIZED_WIRE_2816;
wire	SYNTHESIZED_WIRE_2817;
wire	SYNTHESIZED_WIRE_2818;
wire	SYNTHESIZED_WIRE_2819;
wire	SYNTHESIZED_WIRE_2820;
wire	SYNTHESIZED_WIRE_2821;
wire	SYNTHESIZED_WIRE_2822;
wire	SYNTHESIZED_WIRE_2823;
wire	SYNTHESIZED_WIRE_2824;
wire	SYNTHESIZED_WIRE_2825;
wire	SYNTHESIZED_WIRE_2826;
wire	SYNTHESIZED_WIRE_2827;
wire	SYNTHESIZED_WIRE_2828;
wire	SYNTHESIZED_WIRE_2829;
wire	SYNTHESIZED_WIRE_2830;
wire	SYNTHESIZED_WIRE_2831;
wire	SYNTHESIZED_WIRE_2832;
wire	SYNTHESIZED_WIRE_2833;
wire	SYNTHESIZED_WIRE_2834;
wire	SYNTHESIZED_WIRE_2835;
wire	SYNTHESIZED_WIRE_2836;
wire	SYNTHESIZED_WIRE_2837;
wire	SYNTHESIZED_WIRE_2838;
wire	SYNTHESIZED_WIRE_2839;
wire	SYNTHESIZED_WIRE_2840;
wire	SYNTHESIZED_WIRE_2841;
wire	SYNTHESIZED_WIRE_2842;
wire	SYNTHESIZED_WIRE_2843;
wire	SYNTHESIZED_WIRE_2844;
wire	SYNTHESIZED_WIRE_2845;
wire	SYNTHESIZED_WIRE_2846;
wire	SYNTHESIZED_WIRE_2847;
wire	SYNTHESIZED_WIRE_2848;
wire	SYNTHESIZED_WIRE_2849;
wire	SYNTHESIZED_WIRE_2850;
wire	SYNTHESIZED_WIRE_2851;
wire	SYNTHESIZED_WIRE_2852;
wire	SYNTHESIZED_WIRE_2853;
wire	SYNTHESIZED_WIRE_2854;
wire	SYNTHESIZED_WIRE_2855;
wire	SYNTHESIZED_WIRE_2856;
wire	SYNTHESIZED_WIRE_2857;
wire	SYNTHESIZED_WIRE_2858;
wire	SYNTHESIZED_WIRE_2859;
wire	SYNTHESIZED_WIRE_2860;
wire	SYNTHESIZED_WIRE_2861;
wire	SYNTHESIZED_WIRE_2862;
wire	SYNTHESIZED_WIRE_2863;
wire	SYNTHESIZED_WIRE_2864;
wire	SYNTHESIZED_WIRE_2865;
wire	SYNTHESIZED_WIRE_2866;
wire	SYNTHESIZED_WIRE_2867;
wire	SYNTHESIZED_WIRE_2868;
wire	SYNTHESIZED_WIRE_2869;
wire	SYNTHESIZED_WIRE_2870;
wire	SYNTHESIZED_WIRE_2871;
wire	SYNTHESIZED_WIRE_2872;
wire	SYNTHESIZED_WIRE_2873;
wire	SYNTHESIZED_WIRE_2874;
wire	SYNTHESIZED_WIRE_2875;
wire	SYNTHESIZED_WIRE_2876;
wire	SYNTHESIZED_WIRE_2877;
wire	SYNTHESIZED_WIRE_2878;
wire	SYNTHESIZED_WIRE_2879;
wire	SYNTHESIZED_WIRE_2880;
wire	SYNTHESIZED_WIRE_2881;
wire	SYNTHESIZED_WIRE_2882;
wire	SYNTHESIZED_WIRE_2883;
wire	SYNTHESIZED_WIRE_2884;
wire	SYNTHESIZED_WIRE_2885;
wire	SYNTHESIZED_WIRE_2886;
wire	SYNTHESIZED_WIRE_2887;
wire	SYNTHESIZED_WIRE_2888;
wire	SYNTHESIZED_WIRE_2889;
wire	SYNTHESIZED_WIRE_2890;
wire	SYNTHESIZED_WIRE_2891;
wire	SYNTHESIZED_WIRE_2892;
wire	SYNTHESIZED_WIRE_2893;
wire	SYNTHESIZED_WIRE_2894;
wire	SYNTHESIZED_WIRE_2895;
wire	SYNTHESIZED_WIRE_2896;
wire	SYNTHESIZED_WIRE_2897;
wire	SYNTHESIZED_WIRE_2898;
wire	SYNTHESIZED_WIRE_2899;
wire	SYNTHESIZED_WIRE_2900;
wire	SYNTHESIZED_WIRE_2901;
wire	SYNTHESIZED_WIRE_2902;
wire	SYNTHESIZED_WIRE_2903;
wire	SYNTHESIZED_WIRE_2904;
wire	SYNTHESIZED_WIRE_2905;
wire	SYNTHESIZED_WIRE_2906;
wire	SYNTHESIZED_WIRE_2907;
wire	SYNTHESIZED_WIRE_2908;
wire	SYNTHESIZED_WIRE_2909;
wire	SYNTHESIZED_WIRE_2910;
wire	SYNTHESIZED_WIRE_2911;
wire	SYNTHESIZED_WIRE_2912;
wire	SYNTHESIZED_WIRE_2913;
wire	SYNTHESIZED_WIRE_2914;
wire	SYNTHESIZED_WIRE_2915;
wire	SYNTHESIZED_WIRE_2916;
wire	SYNTHESIZED_WIRE_2917;
wire	SYNTHESIZED_WIRE_2918;
wire	SYNTHESIZED_WIRE_2919;
wire	SYNTHESIZED_WIRE_2920;
wire	SYNTHESIZED_WIRE_2921;
wire	SYNTHESIZED_WIRE_2922;
wire	SYNTHESIZED_WIRE_2923;
wire	SYNTHESIZED_WIRE_2924;
wire	SYNTHESIZED_WIRE_2925;
wire	SYNTHESIZED_WIRE_2926;
wire	SYNTHESIZED_WIRE_2927;
wire	SYNTHESIZED_WIRE_2928;
wire	SYNTHESIZED_WIRE_2929;
wire	SYNTHESIZED_WIRE_2930;
wire	SYNTHESIZED_WIRE_2931;
wire	SYNTHESIZED_WIRE_2932;
wire	SYNTHESIZED_WIRE_2933;
wire	SYNTHESIZED_WIRE_2934;
wire	SYNTHESIZED_WIRE_2935;
wire	SYNTHESIZED_WIRE_2936;
wire	SYNTHESIZED_WIRE_2937;
wire	SYNTHESIZED_WIRE_2938;
wire	SYNTHESIZED_WIRE_2939;
wire	SYNTHESIZED_WIRE_2940;
wire	SYNTHESIZED_WIRE_2941;
wire	SYNTHESIZED_WIRE_2942;
wire	SYNTHESIZED_WIRE_2943;
wire	SYNTHESIZED_WIRE_2944;
wire	SYNTHESIZED_WIRE_2945;
wire	SYNTHESIZED_WIRE_2946;

assign	SYNTHESIZED_WIRE_31 = 1;
assign	SYNTHESIZED_WIRE_674 = 1;





OneBitAdderHalf	b2v_inst1(
	.A(SYNTHESIZED_WIRE_0),
	.B(SYNTHESIZED_WIRE_1),
	.C(SYNTHESIZED_WIRE_1314),
	.S(Z_ALTERA_SYNTHESIZED[31]));


OneBitAdder	b2v_inst100(
	.ci(SYNTHESIZED_WIRE_2),
	.a(SYNTHESIZED_WIRE_3),
	.b(SYNTHESIZED_WIRE_4),
	.co(SYNTHESIZED_WIRE_35),
	.s(SYNTHESIZED_WIRE_1872));


OneBitAdder	b2v_inst1000(
	.ci(SYNTHESIZED_WIRE_5),
	.a(SYNTHESIZED_WIRE_6),
	.b(SYNTHESIZED_WIRE_7),
	.co(SYNTHESIZED_WIRE_8),
	.s(SYNTHESIZED_WIRE_2843));


OneBitAdder	b2v_inst1001(
	.ci(SYNTHESIZED_WIRE_8),
	.a(SYNTHESIZED_WIRE_9),
	.b(SYNTHESIZED_WIRE_10),
	.co(SYNTHESIZED_WIRE_11),
	.s(SYNTHESIZED_WIRE_2846));


OneBitAdder	b2v_inst1002(
	.ci(SYNTHESIZED_WIRE_11),
	.a(SYNTHESIZED_WIRE_12),
	.b(SYNTHESIZED_WIRE_13),
	.co(SYNTHESIZED_WIRE_14),
	.s(SYNTHESIZED_WIRE_2849));


OneBitAdder	b2v_inst1003(
	.ci(SYNTHESIZED_WIRE_14),
	.a(SYNTHESIZED_WIRE_15),
	.b(SYNTHESIZED_WIRE_16),
	.co(SYNTHESIZED_WIRE_17),
	.s(SYNTHESIZED_WIRE_2854));


OneBitAdder	b2v_inst1004(
	.ci(SYNTHESIZED_WIRE_17),
	.a(SYNTHESIZED_WIRE_18),
	.b(SYNTHESIZED_WIRE_19),
	.co(SYNTHESIZED_WIRE_20),
	.s(SYNTHESIZED_WIRE_2857));


OneBitAdder	b2v_inst1005(
	.ci(SYNTHESIZED_WIRE_20),
	.a(SYNTHESIZED_WIRE_21),
	.b(SYNTHESIZED_WIRE_22),
	.co(SYNTHESIZED_WIRE_23),
	.s(SYNTHESIZED_WIRE_2860));


OneBitAdder	b2v_inst1006(
	.ci(SYNTHESIZED_WIRE_23),
	.a(SYNTHESIZED_WIRE_24),
	.b(SYNTHESIZED_WIRE_25),
	.co(SYNTHESIZED_WIRE_26),
	.s(SYNTHESIZED_WIRE_2863));


OneBitAdder	b2v_inst1007(
	.ci(SYNTHESIZED_WIRE_26),
	.a(SYNTHESIZED_WIRE_27),
	.b(SYNTHESIZED_WIRE_28),
	.co(SYNTHESIZED_WIRE_29),
	.s(SYNTHESIZED_WIRE_2866));


OneBitAdder	b2v_inst1008(
	.ci(SYNTHESIZED_WIRE_29),
	.a(SYNTHESIZED_WIRE_30),
	.b(SYNTHESIZED_WIRE_31),
	.co(SYNTHESIZED_WIRE_2872),
	.s(SYNTHESIZED_WIRE_2869));


OneBitAdder	b2v_inst1009(
	.ci(SYNTHESIZED_WIRE_32),
	.a(SYNTHESIZED_WIRE_33),
	.b(SYNTHESIZED_WIRE_34),
	.co(SYNTHESIZED_WIRE_38),
	.s(SYNTHESIZED_WIRE_2824));


OneBitAdder	b2v_inst101(
	.ci(SYNTHESIZED_WIRE_35),
	.a(SYNTHESIZED_WIRE_36),
	.b(SYNTHESIZED_WIRE_37),
	.co(SYNTHESIZED_WIRE_68),
	.s(SYNTHESIZED_WIRE_1904));


OneBitAdder	b2v_inst1010(
	.ci(SYNTHESIZED_WIRE_38),
	.a(SYNTHESIZED_WIRE_39),
	.b(SYNTHESIZED_WIRE_40),
	.co(SYNTHESIZED_WIRE_41),
	.s(SYNTHESIZED_WIRE_2875));


OneBitAdder	b2v_inst1011(
	.ci(SYNTHESIZED_WIRE_41),
	.a(SYNTHESIZED_WIRE_42),
	.b(SYNTHESIZED_WIRE_43),
	.co(SYNTHESIZED_WIRE_44),
	.s(SYNTHESIZED_WIRE_2878));


OneBitAdder	b2v_inst1012(
	.ci(SYNTHESIZED_WIRE_44),
	.a(SYNTHESIZED_WIRE_45),
	.b(SYNTHESIZED_WIRE_46),
	.co(SYNTHESIZED_WIRE_47),
	.s(SYNTHESIZED_WIRE_2881));


OneBitAdder	b2v_inst1013(
	.ci(SYNTHESIZED_WIRE_47),
	.a(SYNTHESIZED_WIRE_48),
	.b(SYNTHESIZED_WIRE_49),
	.co(SYNTHESIZED_WIRE_50),
	.s(SYNTHESIZED_WIRE_2887));


OneBitAdder	b2v_inst1014(
	.ci(SYNTHESIZED_WIRE_50),
	.a(SYNTHESIZED_WIRE_51),
	.b(SYNTHESIZED_WIRE_52),
	.co(SYNTHESIZED_WIRE_53),
	.s(SYNTHESIZED_WIRE_2890));


OneBitAdder	b2v_inst1015(
	.ci(SYNTHESIZED_WIRE_53),
	.a(SYNTHESIZED_WIRE_54),
	.b(SYNTHESIZED_WIRE_55),
	.co(SYNTHESIZED_WIRE_56),
	.s(SYNTHESIZED_WIRE_2893));


OneBitAdder	b2v_inst1016(
	.ci(SYNTHESIZED_WIRE_56),
	.a(SYNTHESIZED_WIRE_57),
	.b(SYNTHESIZED_WIRE_58),
	.co(SYNTHESIZED_WIRE_59),
	.s(SYNTHESIZED_WIRE_2896));


OneBitAdder	b2v_inst1017(
	.ci(SYNTHESIZED_WIRE_59),
	.a(SYNTHESIZED_WIRE_60),
	.b(SYNTHESIZED_WIRE_61),
	.co(SYNTHESIZED_WIRE_62),
	.s(SYNTHESIZED_WIRE_2899));


OneBitAdder	b2v_inst1018(
	.ci(SYNTHESIZED_WIRE_62),
	.a(SYNTHESIZED_WIRE_63),
	.b(SYNTHESIZED_WIRE_64),
	.co(SYNTHESIZED_WIRE_65),
	.s(SYNTHESIZED_WIRE_2902));


OneBitAdder	b2v_inst1019(
	.ci(SYNTHESIZED_WIRE_65),
	.a(SYNTHESIZED_WIRE_66),
	.b(SYNTHESIZED_WIRE_67),
	.co(SYNTHESIZED_WIRE_71),
	.s(SYNTHESIZED_WIRE_2905));


OneBitAdder	b2v_inst102(
	.ci(SYNTHESIZED_WIRE_68),
	.a(SYNTHESIZED_WIRE_69),
	.b(SYNTHESIZED_WIRE_70),
	.co(SYNTHESIZED_WIRE_86),
	.s(SYNTHESIZED_WIRE_1937));


OneBitAdder	b2v_inst1020(
	.ci(SYNTHESIZED_WIRE_71),
	.a(SYNTHESIZED_WIRE_72),
	.b(SYNTHESIZED_WIRE_73),
	.co(SYNTHESIZED_WIRE_74),
	.s(SYNTHESIZED_WIRE_2908));


OneBitAdder	b2v_inst1021(
	.ci(SYNTHESIZED_WIRE_74),
	.a(SYNTHESIZED_WIRE_75),
	.b(SYNTHESIZED_WIRE_76),
	.co(SYNTHESIZED_WIRE_77),
	.s(SYNTHESIZED_WIRE_2911));


OneBitAdder	b2v_inst1022(
	.ci(SYNTHESIZED_WIRE_77),
	.a(SYNTHESIZED_WIRE_78),
	.b(SYNTHESIZED_WIRE_79),
	.co(SYNTHESIZED_WIRE_80),
	.s(SYNTHESIZED_WIRE_2914));


OneBitAdder	b2v_inst1023(
	.ci(SYNTHESIZED_WIRE_80),
	.a(SYNTHESIZED_WIRE_81),
	.b(SYNTHESIZED_WIRE_82),
	.co(SYNTHESIZED_WIRE_83),
	.s(SYNTHESIZED_WIRE_2920));


OneBitAdder	b2v_inst1024(
	.ci(SYNTHESIZED_WIRE_83),
	.a(SYNTHESIZED_WIRE_84),
	.b(SYNTHESIZED_WIRE_85),
	.co(SYNTHESIZED_WIRE_2929),
	.s(SYNTHESIZED_WIRE_2923));

assign	SYNTHESIZED_WIRE_27 = B[1] & A[30];

assign	SYNTHESIZED_WIRE_30 = ~(A[31] & B[1]);

assign	SYNTHESIZED_WIRE_24 = B[1] & A[29];

assign	SYNTHESIZED_WIRE_21 = B[1] & A[28];

assign	SYNTHESIZED_WIRE_18 = B[1] & A[27];


OneBitAdder	b2v_inst103(
	.ci(SYNTHESIZED_WIRE_86),
	.a(SYNTHESIZED_WIRE_87),
	.b(SYNTHESIZED_WIRE_88),
	.co(SYNTHESIZED_WIRE_89),
	.s(SYNTHESIZED_WIRE_1970));

assign	SYNTHESIZED_WIRE_25 = B[0] & A[30];

assign	SYNTHESIZED_WIRE_28 = ~(A[31] & B[0]);

assign	SYNTHESIZED_WIRE_22 = B[0] & A[29];

assign	SYNTHESIZED_WIRE_19 = B[0] & A[28];

assign	SYNTHESIZED_WIRE_15 = B[1] & A[26];

assign	SYNTHESIZED_WIRE_12 = B[1] & A[25];

assign	SYNTHESIZED_WIRE_9 = B[1] & A[24];

assign	SYNTHESIZED_WIRE_6 = B[1] & A[23];

assign	SYNTHESIZED_WIRE_2945 = B[1] & A[22];

assign	SYNTHESIZED_WIRE_2942 = B[1] & A[21];


OneBitAdder	b2v_inst104(
	.ci(SYNTHESIZED_WIRE_89),
	.a(SYNTHESIZED_WIRE_90),
	.b(SYNTHESIZED_WIRE_91),
	.co(SYNTHESIZED_WIRE_92),
	.s(SYNTHESIZED_WIRE_2002));

assign	SYNTHESIZED_WIRE_2939 = B[1] & A[20];

assign	SYNTHESIZED_WIRE_2936 = B[1] & A[19];

assign	SYNTHESIZED_WIRE_2933 = B[1] & A[18];

assign	SYNTHESIZED_WIRE_2930 = B[1] & A[17];

assign	SYNTHESIZED_WIRE_84 = B[1] & A[16];

assign	SYNTHESIZED_WIRE_81 = B[1] & A[15];

assign	SYNTHESIZED_WIRE_78 = B[1] & A[14];

assign	SYNTHESIZED_WIRE_75 = B[1] & A[13];

assign	SYNTHESIZED_WIRE_72 = B[1] & A[12];

assign	SYNTHESIZED_WIRE_66 = B[1] & A[11];


OneBitAdder	b2v_inst105(
	.ci(SYNTHESIZED_WIRE_92),
	.a(SYNTHESIZED_WIRE_93),
	.b(SYNTHESIZED_WIRE_94),
	.co(SYNTHESIZED_WIRE_95),
	.s(SYNTHESIZED_WIRE_2035));

assign	SYNTHESIZED_WIRE_63 = B[1] & A[10];

assign	SYNTHESIZED_WIRE_60 = B[1] & A[9];

assign	SYNTHESIZED_WIRE_57 = B[1] & A[8];

assign	SYNTHESIZED_WIRE_54 = B[1] & A[7];

assign	SYNTHESIZED_WIRE_51 = B[1] & A[6];

assign	SYNTHESIZED_WIRE_48 = B[1] & A[5];

assign	SYNTHESIZED_WIRE_45 = B[1] & A[4];

assign	SYNTHESIZED_WIRE_42 = B[1] & A[3];

assign	SYNTHESIZED_WIRE_39 = B[1] & A[2];

assign	SYNTHESIZED_WIRE_33 = B[1] & A[1];


OneBitAdder	b2v_inst106(
	.ci(SYNTHESIZED_WIRE_95),
	.a(SYNTHESIZED_WIRE_96),
	.b(SYNTHESIZED_WIRE_97),
	.co(SYNTHESIZED_WIRE_98),
	.s(SYNTHESIZED_WIRE_2068));

assign	SYNTHESIZED_WIRE_2928 = B[1] & A[0];

assign	SYNTHESIZED_WIRE_16 = B[0] & A[27];

assign	SYNTHESIZED_WIRE_13 = B[0] & A[26];

assign	SYNTHESIZED_WIRE_10 = B[0] & A[25];

assign	SYNTHESIZED_WIRE_7 = B[0] & A[24];

assign	SYNTHESIZED_WIRE_2946 = B[0] & A[23];

assign	SYNTHESIZED_WIRE_2943 = B[0] & A[22];

assign	SYNTHESIZED_WIRE_2940 = B[0] & A[21];

assign	SYNTHESIZED_WIRE_2937 = B[0] & A[20];

assign	SYNTHESIZED_WIRE_2934 = B[0] & A[19];


OneBitAdder	b2v_inst107(
	.ci(SYNTHESIZED_WIRE_98),
	.a(SYNTHESIZED_WIRE_99),
	.b(SYNTHESIZED_WIRE_100),
	.co(SYNTHESIZED_WIRE_101),
	.s(SYNTHESIZED_WIRE_2100));

assign	SYNTHESIZED_WIRE_2931 = B[0] & A[18];

assign	SYNTHESIZED_WIRE_85 = B[0] & A[17];

assign	SYNTHESIZED_WIRE_82 = B[0] & A[16];

assign	SYNTHESIZED_WIRE_79 = B[0] & A[15];

assign	SYNTHESIZED_WIRE_76 = B[0] & A[14];

assign	SYNTHESIZED_WIRE_73 = B[0] & A[13];

assign	SYNTHESIZED_WIRE_67 = B[0] & A[12];

assign	SYNTHESIZED_WIRE_64 = B[0] & A[11];

assign	SYNTHESIZED_WIRE_61 = B[0] & A[10];

assign	SYNTHESIZED_WIRE_58 = B[0] & A[9];


OneBitAdder	b2v_inst108(
	.ci(SYNTHESIZED_WIRE_101),
	.a(SYNTHESIZED_WIRE_102),
	.b(SYNTHESIZED_WIRE_103),
	.co(SYNTHESIZED_WIRE_104),
	.s(SYNTHESIZED_WIRE_2133));

assign	SYNTHESIZED_WIRE_55 = B[0] & A[8];

assign	SYNTHESIZED_WIRE_52 = B[0] & A[7];

assign	SYNTHESIZED_WIRE_49 = B[0] & A[6];

assign	SYNTHESIZED_WIRE_46 = B[0] & A[5];

assign	SYNTHESIZED_WIRE_43 = B[0] & A[4];

assign	SYNTHESIZED_WIRE_40 = B[0] & A[3];

assign	SYNTHESIZED_WIRE_34 = B[0] & A[2];

assign	SYNTHESIZED_WIRE_2927 = B[0] & A[1];

assign	Z_ALTERA_SYNTHESIZED[0] = B[0] & A[0];

assign	SYNTHESIZED_WIRE_2868 = B[2] & A[30];


OneBitAdder	b2v_inst109(
	.ci(SYNTHESIZED_WIRE_104),
	.a(SYNTHESIZED_WIRE_105),
	.b(SYNTHESIZED_WIRE_106),
	.co(SYNTHESIZED_WIRE_107),
	.s(SYNTHESIZED_WIRE_2166));

assign	SYNTHESIZED_WIRE_2871 = ~(A[31] & B[2]);

assign	SYNTHESIZED_WIRE_2865 = B[2] & A[29];

assign	SYNTHESIZED_WIRE_2862 = B[2] & A[28];

assign	SYNTHESIZED_WIRE_2859 = B[2] & A[27];

assign	SYNTHESIZED_WIRE_2856 = B[2] & A[26];

assign	SYNTHESIZED_WIRE_2853 = B[2] & A[25];

assign	SYNTHESIZED_WIRE_2848 = B[2] & A[24];

assign	SYNTHESIZED_WIRE_2845 = B[2] & A[23];

assign	SYNTHESIZED_WIRE_2842 = B[2] & A[22];

assign	SYNTHESIZED_WIRE_2839 = B[2] & A[21];


OneBitAdder	b2v_inst110(
	.ci(SYNTHESIZED_WIRE_107),
	.a(SYNTHESIZED_WIRE_108),
	.b(SYNTHESIZED_WIRE_109),
	.co(SYNTHESIZED_WIRE_110),
	.s(SYNTHESIZED_WIRE_2198));

assign	SYNTHESIZED_WIRE_2836 = B[2] & A[20];

assign	SYNTHESIZED_WIRE_2833 = B[2] & A[19];

assign	SYNTHESIZED_WIRE_2830 = B[2] & A[18];

assign	SYNTHESIZED_WIRE_2827 = B[2] & A[17];

assign	SYNTHESIZED_WIRE_2925 = B[2] & A[16];

assign	SYNTHESIZED_WIRE_2922 = B[2] & A[15];

assign	SYNTHESIZED_WIRE_2919 = B[2] & A[14];

assign	SYNTHESIZED_WIRE_2913 = B[2] & A[13];

assign	SYNTHESIZED_WIRE_2910 = B[2] & A[12];

assign	SYNTHESIZED_WIRE_2907 = B[2] & A[11];


OneBitAdder	b2v_inst111(
	.ci(SYNTHESIZED_WIRE_110),
	.a(SYNTHESIZED_WIRE_111),
	.b(SYNTHESIZED_WIRE_112),
	.co(SYNTHESIZED_WIRE_113),
	.s(SYNTHESIZED_WIRE_2231));

assign	SYNTHESIZED_WIRE_2904 = B[2] & A[10];

assign	SYNTHESIZED_WIRE_2901 = B[2] & A[9];

assign	SYNTHESIZED_WIRE_2898 = B[2] & A[8];

assign	SYNTHESIZED_WIRE_2895 = B[2] & A[7];

assign	SYNTHESIZED_WIRE_2892 = B[2] & A[6];

assign	SYNTHESIZED_WIRE_2889 = B[2] & A[5];

assign	SYNTHESIZED_WIRE_2886 = B[2] & A[4];

assign	SYNTHESIZED_WIRE_2880 = B[2] & A[3];

assign	SYNTHESIZED_WIRE_2877 = B[2] & A[2];

assign	SYNTHESIZED_WIRE_2874 = B[2] & A[1];


OneBitAdder	b2v_inst112(
	.ci(SYNTHESIZED_WIRE_113),
	.a(SYNTHESIZED_WIRE_114),
	.b(SYNTHESIZED_WIRE_115),
	.co(SYNTHESIZED_WIRE_2297),
	.s(SYNTHESIZED_WIRE_2264));

assign	SYNTHESIZED_WIRE_2825 = B[2] & A[0];

assign	SYNTHESIZED_WIRE_2765 = B[3] & A[30];

assign	SYNTHESIZED_WIRE_2768 = ~(A[31] & B[3]);

assign	SYNTHESIZED_WIRE_2762 = B[3] & A[29];

assign	SYNTHESIZED_WIRE_2759 = B[3] & A[28];

assign	SYNTHESIZED_WIRE_2756 = B[3] & A[27];

assign	SYNTHESIZED_WIRE_2750 = B[3] & A[26];

assign	SYNTHESIZED_WIRE_2747 = B[3] & A[25];

assign	SYNTHESIZED_WIRE_2744 = B[3] & A[24];

assign	SYNTHESIZED_WIRE_2741 = B[3] & A[23];


OneBitAdder	b2v_inst113(
	.ci(SYNTHESIZED_WIRE_116),
	.a(SYNTHESIZED_WIRE_117),
	.b(SYNTHESIZED_WIRE_118),
	.co(SYNTHESIZED_WIRE_119),
	.s(SYNTHESIZED_WIRE_374));

assign	SYNTHESIZED_WIRE_2738 = B[3] & A[22];

assign	SYNTHESIZED_WIRE_2735 = B[3] & A[21];

assign	SYNTHESIZED_WIRE_2732 = B[3] & A[20];

assign	SYNTHESIZED_WIRE_2729 = B[3] & A[19];

assign	SYNTHESIZED_WIRE_2726 = B[3] & A[18];

assign	SYNTHESIZED_WIRE_2723 = B[3] & A[17];

assign	SYNTHESIZED_WIRE_2822 = B[3] & A[16];

assign	SYNTHESIZED_WIRE_2816 = B[3] & A[15];

assign	SYNTHESIZED_WIRE_2813 = B[3] & A[14];

assign	SYNTHESIZED_WIRE_2810 = B[3] & A[13];


OneBitAdder	b2v_inst114(
	.ci(SYNTHESIZED_WIRE_119),
	.a(SYNTHESIZED_WIRE_120),
	.b(SYNTHESIZED_WIRE_121),
	.co(SYNTHESIZED_WIRE_122),
	.s(SYNTHESIZED_WIRE_2329));

assign	SYNTHESIZED_WIRE_2807 = B[3] & A[12];

assign	SYNTHESIZED_WIRE_2804 = B[3] & A[11];

assign	SYNTHESIZED_WIRE_2801 = B[3] & A[10];

assign	SYNTHESIZED_WIRE_2798 = B[3] & A[9];

assign	SYNTHESIZED_WIRE_2795 = B[3] & A[8];

assign	SYNTHESIZED_WIRE_2792 = B[3] & A[7];

assign	SYNTHESIZED_WIRE_2789 = B[3] & A[6];

assign	SYNTHESIZED_WIRE_2783 = B[3] & A[5];

assign	SYNTHESIZED_WIRE_2780 = B[3] & A[4];

assign	SYNTHESIZED_WIRE_2777 = B[3] & A[3];


OneBitAdder	b2v_inst115(
	.ci(SYNTHESIZED_WIRE_122),
	.a(SYNTHESIZED_WIRE_123),
	.b(SYNTHESIZED_WIRE_124),
	.co(SYNTHESIZED_WIRE_125),
	.s(SYNTHESIZED_WIRE_2362));

assign	SYNTHESIZED_WIRE_2774 = B[3] & A[2];

assign	SYNTHESIZED_WIRE_2771 = B[3] & A[1];

assign	SYNTHESIZED_WIRE_2718 = B[3] & A[0];

assign	SYNTHESIZED_WIRE_2661 = B[4] & A[30];

assign	SYNTHESIZED_WIRE_2664 = ~(A[31] & B[4]);

assign	SYNTHESIZED_WIRE_2658 = B[4] & A[29];

assign	SYNTHESIZED_WIRE_2652 = B[4] & A[28];

assign	SYNTHESIZED_WIRE_2649 = B[4] & A[27];

assign	SYNTHESIZED_WIRE_2646 = B[4] & A[26];

assign	SYNTHESIZED_WIRE_2643 = B[4] & A[25];


OneBitAdder	b2v_inst116(
	.ci(SYNTHESIZED_WIRE_125),
	.a(SYNTHESIZED_WIRE_126),
	.b(SYNTHESIZED_WIRE_127),
	.co(SYNTHESIZED_WIRE_128),
	.s(SYNTHESIZED_WIRE_2395));

assign	SYNTHESIZED_WIRE_2640 = B[4] & A[24];

assign	SYNTHESIZED_WIRE_2637 = B[4] & A[23];

assign	SYNTHESIZED_WIRE_2634 = B[4] & A[22];

assign	SYNTHESIZED_WIRE_2631 = B[4] & A[21];

assign	SYNTHESIZED_WIRE_2628 = B[4] & A[20];

assign	SYNTHESIZED_WIRE_2625 = B[4] & A[19];

assign	SYNTHESIZED_WIRE_2619 = B[4] & A[18];

assign	SYNTHESIZED_WIRE_2616 = B[4] & A[17];

assign	SYNTHESIZED_WIRE_2715 = B[4] & A[16];

assign	SYNTHESIZED_WIRE_2712 = B[4] & A[15];


OneBitAdder	b2v_inst117(
	.ci(SYNTHESIZED_WIRE_128),
	.a(SYNTHESIZED_WIRE_129),
	.b(SYNTHESIZED_WIRE_130),
	.co(SYNTHESIZED_WIRE_131),
	.s(SYNTHESIZED_WIRE_2427));

assign	SYNTHESIZED_WIRE_2709 = B[4] & A[14];

assign	SYNTHESIZED_WIRE_2706 = B[4] & A[13];

assign	SYNTHESIZED_WIRE_2703 = B[4] & A[12];

assign	SYNTHESIZED_WIRE_2700 = B[4] & A[11];

assign	SYNTHESIZED_WIRE_2697 = B[4] & A[10];

assign	SYNTHESIZED_WIRE_2694 = B[4] & A[9];

assign	SYNTHESIZED_WIRE_2691 = B[4] & A[8];

assign	SYNTHESIZED_WIRE_2685 = B[4] & A[7];

assign	SYNTHESIZED_WIRE_2682 = B[4] & A[6];

assign	SYNTHESIZED_WIRE_2679 = B[4] & A[5];


OneBitAdder	b2v_inst118(
	.ci(SYNTHESIZED_WIRE_131),
	.a(SYNTHESIZED_WIRE_132),
	.b(SYNTHESIZED_WIRE_133),
	.co(SYNTHESIZED_WIRE_134),
	.s(SYNTHESIZED_WIRE_2460));

assign	SYNTHESIZED_WIRE_2676 = B[4] & A[4];

assign	SYNTHESIZED_WIRE_2673 = B[4] & A[3];

assign	SYNTHESIZED_WIRE_2670 = B[4] & A[2];

assign	SYNTHESIZED_WIRE_2667 = B[4] & A[1];

assign	SYNTHESIZED_WIRE_2614 = B[4] & A[0];

assign	SYNTHESIZED_WIRE_2554 = B[5] & A[30];

assign	SYNTHESIZED_WIRE_2560 = ~(A[31] & B[5]);

assign	SYNTHESIZED_WIRE_2551 = B[5] & A[29];

assign	SYNTHESIZED_WIRE_2548 = B[5] & A[28];

assign	SYNTHESIZED_WIRE_2545 = B[5] & A[27];


OneBitAdder	b2v_inst119(
	.ci(SYNTHESIZED_WIRE_134),
	.a(SYNTHESIZED_WIRE_135),
	.b(SYNTHESIZED_WIRE_136),
	.co(SYNTHESIZED_WIRE_137),
	.s(SYNTHESIZED_WIRE_2493));

assign	SYNTHESIZED_WIRE_2542 = B[5] & A[26];

assign	SYNTHESIZED_WIRE_2539 = B[5] & A[25];

assign	SYNTHESIZED_WIRE_2536 = B[5] & A[24];

assign	SYNTHESIZED_WIRE_2533 = B[5] & A[23];

assign	SYNTHESIZED_WIRE_2530 = B[5] & A[22];

assign	SYNTHESIZED_WIRE_2527 = B[5] & A[21];

assign	SYNTHESIZED_WIRE_2521 = B[5] & A[20];

assign	SYNTHESIZED_WIRE_2518 = B[5] & A[19];

assign	SYNTHESIZED_WIRE_2515 = B[5] & A[18];

assign	SYNTHESIZED_WIRE_2512 = B[5] & A[17];


OneBitAdder	b2v_inst120(
	.ci(SYNTHESIZED_WIRE_137),
	.a(SYNTHESIZED_WIRE_138),
	.b(SYNTHESIZED_WIRE_139),
	.co(SYNTHESIZED_WIRE_140),
	.s(SYNTHESIZED_WIRE_2525));

assign	SYNTHESIZED_WIRE_2611 = B[5] & A[16];

assign	SYNTHESIZED_WIRE_2608 = B[5] & A[15];

assign	SYNTHESIZED_WIRE_2605 = B[5] & A[14];

assign	SYNTHESIZED_WIRE_2602 = B[5] & A[13];

assign	SYNTHESIZED_WIRE_2599 = B[5] & A[12];

assign	SYNTHESIZED_WIRE_2596 = B[5] & A[11];

assign	SYNTHESIZED_WIRE_2593 = B[5] & A[10];

assign	SYNTHESIZED_WIRE_2587 = B[5] & A[9];

assign	SYNTHESIZED_WIRE_2584 = B[5] & A[8];

assign	SYNTHESIZED_WIRE_2581 = B[5] & A[7];


OneBitAdder	b2v_inst121(
	.ci(SYNTHESIZED_WIRE_140),
	.a(SYNTHESIZED_WIRE_141),
	.b(SYNTHESIZED_WIRE_142),
	.co(SYNTHESIZED_WIRE_143),
	.s(SYNTHESIZED_WIRE_2558));

assign	SYNTHESIZED_WIRE_2578 = B[5] & A[6];

assign	SYNTHESIZED_WIRE_2575 = B[5] & A[5];

assign	SYNTHESIZED_WIRE_2572 = B[5] & A[4];

assign	SYNTHESIZED_WIRE_2569 = B[5] & A[3];

assign	SYNTHESIZED_WIRE_2566 = B[5] & A[2];

assign	SYNTHESIZED_WIRE_2563 = B[5] & A[1];

assign	SYNTHESIZED_WIRE_2510 = B[5] & A[0];

assign	SYNTHESIZED_WIRE_2450 = B[6] & A[30];

assign	SYNTHESIZED_WIRE_2453 = ~(A[31] & B[6]);

assign	SYNTHESIZED_WIRE_2447 = B[6] & A[29];


OneBitAdder	b2v_inst122(
	.ci(SYNTHESIZED_WIRE_143),
	.a(SYNTHESIZED_WIRE_144),
	.b(SYNTHESIZED_WIRE_145),
	.co(SYNTHESIZED_WIRE_146),
	.s(SYNTHESIZED_WIRE_2591));

assign	SYNTHESIZED_WIRE_2444 = B[6] & A[28];

assign	SYNTHESIZED_WIRE_2441 = B[6] & A[27];

assign	SYNTHESIZED_WIRE_2438 = B[6] & A[26];

assign	SYNTHESIZED_WIRE_2435 = B[6] & A[25];

assign	SYNTHESIZED_WIRE_2432 = B[6] & A[24];

assign	SYNTHESIZED_WIRE_2429 = B[6] & A[23];

assign	SYNTHESIZED_WIRE_2423 = B[6] & A[22];

assign	SYNTHESIZED_WIRE_2420 = B[6] & A[21];

assign	SYNTHESIZED_WIRE_2417 = B[6] & A[20];

assign	SYNTHESIZED_WIRE_2414 = B[6] & A[19];


OneBitAdder	b2v_inst123(
	.ci(SYNTHESIZED_WIRE_146),
	.a(SYNTHESIZED_WIRE_147),
	.b(SYNTHESIZED_WIRE_148),
	.co(SYNTHESIZED_WIRE_149),
	.s(SYNTHESIZED_WIRE_2623));

assign	SYNTHESIZED_WIRE_2411 = B[6] & A[18];

assign	SYNTHESIZED_WIRE_2408 = B[6] & A[17];

assign	SYNTHESIZED_WIRE_2507 = B[6] & A[16];

assign	SYNTHESIZED_WIRE_2504 = B[6] & A[15];

assign	SYNTHESIZED_WIRE_2501 = B[6] & A[14];

assign	SYNTHESIZED_WIRE_2498 = B[6] & A[13];

assign	SYNTHESIZED_WIRE_2495 = B[6] & A[12];

assign	SYNTHESIZED_WIRE_2489 = B[6] & A[11];

assign	SYNTHESIZED_WIRE_2486 = B[6] & A[10];

assign	SYNTHESIZED_WIRE_2483 = B[6] & A[9];


OneBitAdder	b2v_inst124(
	.ci(SYNTHESIZED_WIRE_149),
	.a(SYNTHESIZED_WIRE_150),
	.b(SYNTHESIZED_WIRE_151),
	.co(SYNTHESIZED_WIRE_152),
	.s(SYNTHESIZED_WIRE_2656));

assign	SYNTHESIZED_WIRE_2480 = B[6] & A[8];

assign	SYNTHESIZED_WIRE_2477 = B[6] & A[7];

assign	SYNTHESIZED_WIRE_2474 = B[6] & A[6];

assign	SYNTHESIZED_WIRE_2471 = B[6] & A[5];

assign	SYNTHESIZED_WIRE_2468 = B[6] & A[4];

assign	SYNTHESIZED_WIRE_2465 = B[6] & A[3];

assign	SYNTHESIZED_WIRE_2462 = B[6] & A[2];

assign	SYNTHESIZED_WIRE_2456 = B[6] & A[1];

assign	SYNTHESIZED_WIRE_2406 = B[6] & A[0];

assign	SYNTHESIZED_WIRE_2346 = B[7] & A[30];


OneBitAdder	b2v_inst125(
	.ci(SYNTHESIZED_WIRE_152),
	.a(SYNTHESIZED_WIRE_153),
	.b(SYNTHESIZED_WIRE_154),
	.co(SYNTHESIZED_WIRE_155),
	.s(SYNTHESIZED_WIRE_2689));

assign	SYNTHESIZED_WIRE_2349 = ~(A[31] & B[7]);

assign	SYNTHESIZED_WIRE_2343 = B[7] & A[29];

assign	SYNTHESIZED_WIRE_2340 = B[7] & A[28];

assign	SYNTHESIZED_WIRE_2337 = B[7] & A[27];

assign	SYNTHESIZED_WIRE_2334 = B[7] & A[26];

assign	SYNTHESIZED_WIRE_2331 = B[7] & A[25];

assign	SYNTHESIZED_WIRE_2325 = B[7] & A[24];

assign	SYNTHESIZED_WIRE_2322 = B[7] & A[23];

assign	SYNTHESIZED_WIRE_2319 = B[7] & A[22];

assign	SYNTHESIZED_WIRE_2316 = B[7] & A[21];


OneBitAdder	b2v_inst126(
	.ci(SYNTHESIZED_WIRE_155),
	.a(SYNTHESIZED_WIRE_156),
	.b(SYNTHESIZED_WIRE_157),
	.co(SYNTHESIZED_WIRE_158),
	.s(SYNTHESIZED_WIRE_2721));

assign	SYNTHESIZED_WIRE_2313 = B[7] & A[20];

assign	SYNTHESIZED_WIRE_2310 = B[7] & A[19];

assign	SYNTHESIZED_WIRE_2307 = B[7] & A[18];

assign	SYNTHESIZED_WIRE_2304 = B[7] & A[17];

assign	SYNTHESIZED_WIRE_2403 = B[7] & A[16];

assign	SYNTHESIZED_WIRE_2400 = B[7] & A[15];

assign	SYNTHESIZED_WIRE_2397 = B[7] & A[14];

assign	SYNTHESIZED_WIRE_2391 = B[7] & A[13];

assign	SYNTHESIZED_WIRE_2388 = B[7] & A[12];

assign	SYNTHESIZED_WIRE_2385 = B[7] & A[11];


OneBitAdder	b2v_inst127(
	.ci(SYNTHESIZED_WIRE_158),
	.a(SYNTHESIZED_WIRE_159),
	.b(SYNTHESIZED_WIRE_160),
	.co(SYNTHESIZED_WIRE_161),
	.s(SYNTHESIZED_WIRE_2754));

assign	SYNTHESIZED_WIRE_2382 = B[7] & A[10];

assign	SYNTHESIZED_WIRE_2379 = B[7] & A[9];

assign	SYNTHESIZED_WIRE_2376 = B[7] & A[8];

assign	SYNTHESIZED_WIRE_2373 = B[7] & A[7];

assign	SYNTHESIZED_WIRE_2370 = B[7] & A[6];

assign	SYNTHESIZED_WIRE_2367 = B[7] & A[5];

assign	SYNTHESIZED_WIRE_2364 = B[7] & A[4];

assign	SYNTHESIZED_WIRE_2358 = B[7] & A[3];

assign	SYNTHESIZED_WIRE_2355 = B[7] & A[2];

assign	SYNTHESIZED_WIRE_2352 = B[7] & A[1];


OneBitAdder	b2v_inst128(
	.ci(SYNTHESIZED_WIRE_161),
	.a(SYNTHESIZED_WIRE_162),
	.b(SYNTHESIZED_WIRE_163),
	.co(SYNTHESIZED_WIRE_2882),
	.s(SYNTHESIZED_WIRE_2787));

assign	SYNTHESIZED_WIRE_2302 = B[7] & A[0];

assign	SYNTHESIZED_WIRE_2242 = B[8] & A[30];

assign	SYNTHESIZED_WIRE_2245 = ~(A[31] & B[8]);

assign	SYNTHESIZED_WIRE_2239 = B[8] & A[29];

assign	SYNTHESIZED_WIRE_2236 = B[8] & A[28];

assign	SYNTHESIZED_WIRE_2233 = B[8] & A[27];

assign	SYNTHESIZED_WIRE_2227 = B[8] & A[26];

assign	SYNTHESIZED_WIRE_2224 = B[8] & A[25];

assign	SYNTHESIZED_WIRE_2221 = B[8] & A[24];

assign	SYNTHESIZED_WIRE_2218 = B[8] & A[23];


OneBitAdderHalf	b2v_inst129(
	.A(SYNTHESIZED_WIRE_164),
	.B(SYNTHESIZED_WIRE_165),
	.C(SYNTHESIZED_WIRE_211),
	.S(Z_ALTERA_SYNTHESIZED[28]));

assign	SYNTHESIZED_WIRE_2215 = B[8] & A[22];

assign	SYNTHESIZED_WIRE_2212 = B[8] & A[21];

assign	SYNTHESIZED_WIRE_2209 = B[8] & A[20];

assign	SYNTHESIZED_WIRE_2206 = B[8] & A[19];

assign	SYNTHESIZED_WIRE_2203 = B[8] & A[18];

assign	SYNTHESIZED_WIRE_2200 = B[8] & A[17];

assign	SYNTHESIZED_WIRE_2299 = B[8] & A[16];

assign	SYNTHESIZED_WIRE_2293 = B[8] & A[15];

assign	SYNTHESIZED_WIRE_2290 = B[8] & A[14];

assign	SYNTHESIZED_WIRE_2287 = B[8] & A[13];


OneBitAdder	b2v_inst130(
	.ci(SYNTHESIZED_WIRE_166),
	.a(SYNTHESIZED_WIRE_167),
	.b(SYNTHESIZED_WIRE_168),
	.co(SYNTHESIZED_WIRE_169),
	.s(SYNTHESIZED_WIRE_163));

assign	SYNTHESIZED_WIRE_2284 = B[8] & A[12];

assign	SYNTHESIZED_WIRE_2281 = B[8] & A[11];

assign	SYNTHESIZED_WIRE_2278 = B[8] & A[10];

assign	SYNTHESIZED_WIRE_2275 = B[8] & A[9];

assign	SYNTHESIZED_WIRE_2272 = B[8] & A[8];

assign	SYNTHESIZED_WIRE_2269 = B[8] & A[7];

assign	SYNTHESIZED_WIRE_2266 = B[8] & A[6];

assign	SYNTHESIZED_WIRE_2260 = B[8] & A[5];

assign	SYNTHESIZED_WIRE_2257 = B[8] & A[4];

assign	SYNTHESIZED_WIRE_2254 = B[8] & A[3];


OneBitAdder	b2v_inst131(
	.ci(SYNTHESIZED_WIRE_169),
	.a(SYNTHESIZED_WIRE_170),
	.b(SYNTHESIZED_WIRE_171),
	.co(SYNTHESIZED_WIRE_172),
	.s(SYNTHESIZED_WIRE_2884));

assign	SYNTHESIZED_WIRE_2251 = B[8] & A[2];

assign	SYNTHESIZED_WIRE_2248 = B[8] & A[1];

assign	SYNTHESIZED_WIRE_2195 = B[8] & A[0];

assign	SYNTHESIZED_WIRE_2138 = B[9] & A[30];

assign	SYNTHESIZED_WIRE_2141 = ~(A[31] & B[9]);

assign	SYNTHESIZED_WIRE_2135 = B[9] & A[29];

assign	SYNTHESIZED_WIRE_2129 = B[9] & A[28];

assign	SYNTHESIZED_WIRE_2126 = B[9] & A[27];

assign	SYNTHESIZED_WIRE_2123 = B[9] & A[26];

assign	SYNTHESIZED_WIRE_2120 = B[9] & A[25];


OneBitAdder	b2v_inst132(
	.ci(SYNTHESIZED_WIRE_172),
	.a(SYNTHESIZED_WIRE_173),
	.b(SYNTHESIZED_WIRE_174),
	.co(SYNTHESIZED_WIRE_175),
	.s(SYNTHESIZED_WIRE_2917));

assign	SYNTHESIZED_WIRE_2117 = B[9] & A[24];

assign	SYNTHESIZED_WIRE_2114 = B[9] & A[23];

assign	SYNTHESIZED_WIRE_2111 = B[9] & A[22];

assign	SYNTHESIZED_WIRE_2108 = B[9] & A[21];

assign	SYNTHESIZED_WIRE_2105 = B[9] & A[20];

assign	SYNTHESIZED_WIRE_2102 = B[9] & A[19];

assign	SYNTHESIZED_WIRE_2096 = B[9] & A[18];

assign	SYNTHESIZED_WIRE_2093 = B[9] & A[17];

assign	SYNTHESIZED_WIRE_2192 = B[9] & A[16];

assign	SYNTHESIZED_WIRE_2189 = B[9] & A[15];


OneBitAdder	b2v_inst133(
	.ci(SYNTHESIZED_WIRE_175),
	.a(SYNTHESIZED_WIRE_176),
	.b(SYNTHESIZED_WIRE_177),
	.co(SYNTHESIZED_WIRE_178),
	.s(SYNTHESIZED_WIRE_4));

assign	SYNTHESIZED_WIRE_2186 = B[9] & A[14];

assign	SYNTHESIZED_WIRE_2183 = B[9] & A[13];

assign	SYNTHESIZED_WIRE_2180 = B[9] & A[12];

assign	SYNTHESIZED_WIRE_2177 = B[9] & A[11];

assign	SYNTHESIZED_WIRE_2174 = B[9] & A[10];

assign	SYNTHESIZED_WIRE_2171 = B[9] & A[9];

assign	SYNTHESIZED_WIRE_2168 = B[9] & A[8];

assign	SYNTHESIZED_WIRE_2162 = B[9] & A[7];

assign	SYNTHESIZED_WIRE_2159 = B[9] & A[6];

assign	SYNTHESIZED_WIRE_2156 = B[9] & A[5];


OneBitAdder	b2v_inst134(
	.ci(SYNTHESIZED_WIRE_178),
	.a(SYNTHESIZED_WIRE_179),
	.b(SYNTHESIZED_WIRE_180),
	.co(SYNTHESIZED_WIRE_181),
	.s(SYNTHESIZED_WIRE_37));

assign	SYNTHESIZED_WIRE_2153 = B[9] & A[4];

assign	SYNTHESIZED_WIRE_2150 = B[9] & A[3];

assign	SYNTHESIZED_WIRE_2147 = B[9] & A[2];

assign	SYNTHESIZED_WIRE_2144 = B[9] & A[1];

assign	SYNTHESIZED_WIRE_2091 = B[9] & A[0];

assign	SYNTHESIZED_WIRE_2031 = B[10] & A[30];

assign	SYNTHESIZED_WIRE_2037 = ~(A[31] & B[10]);

assign	SYNTHESIZED_WIRE_2028 = B[10] & A[29];

assign	SYNTHESIZED_WIRE_2025 = B[10] & A[28];

assign	SYNTHESIZED_WIRE_2022 = B[10] & A[27];


OneBitAdder	b2v_inst135(
	.ci(SYNTHESIZED_WIRE_181),
	.a(SYNTHESIZED_WIRE_182),
	.b(SYNTHESIZED_WIRE_183),
	.co(SYNTHESIZED_WIRE_184),
	.s(SYNTHESIZED_WIRE_70));

assign	SYNTHESIZED_WIRE_2019 = B[10] & A[26];

assign	SYNTHESIZED_WIRE_2016 = B[10] & A[25];

assign	SYNTHESIZED_WIRE_2013 = B[10] & A[24];

assign	SYNTHESIZED_WIRE_2010 = B[10] & A[23];

assign	SYNTHESIZED_WIRE_2007 = B[10] & A[22];

assign	SYNTHESIZED_WIRE_2004 = B[10] & A[21];

assign	SYNTHESIZED_WIRE_1998 = B[10] & A[20];

assign	SYNTHESIZED_WIRE_1995 = B[10] & A[19];

assign	SYNTHESIZED_WIRE_1992 = B[10] & A[18];

assign	SYNTHESIZED_WIRE_1989 = B[10] & A[17];


OneBitAdder	b2v_inst136(
	.ci(SYNTHESIZED_WIRE_184),
	.a(SYNTHESIZED_WIRE_185),
	.b(SYNTHESIZED_WIRE_186),
	.co(SYNTHESIZED_WIRE_187),
	.s(SYNTHESIZED_WIRE_88));

assign	SYNTHESIZED_WIRE_2088 = B[10] & A[16];

assign	SYNTHESIZED_WIRE_2085 = B[10] & A[15];

assign	SYNTHESIZED_WIRE_2082 = B[10] & A[14];

assign	SYNTHESIZED_WIRE_2079 = B[10] & A[13];

assign	SYNTHESIZED_WIRE_2076 = B[10] & A[12];

assign	SYNTHESIZED_WIRE_2073 = B[10] & A[11];

assign	SYNTHESIZED_WIRE_2070 = B[10] & A[10];

assign	SYNTHESIZED_WIRE_2064 = B[10] & A[9];

assign	SYNTHESIZED_WIRE_2061 = B[10] & A[8];

assign	SYNTHESIZED_WIRE_2058 = B[10] & A[7];


OneBitAdder	b2v_inst137(
	.ci(SYNTHESIZED_WIRE_187),
	.a(SYNTHESIZED_WIRE_188),
	.b(SYNTHESIZED_WIRE_189),
	.co(SYNTHESIZED_WIRE_190),
	.s(SYNTHESIZED_WIRE_91));

assign	SYNTHESIZED_WIRE_2055 = B[10] & A[6];

assign	SYNTHESIZED_WIRE_2052 = B[10] & A[5];

assign	SYNTHESIZED_WIRE_2049 = B[10] & A[4];

assign	SYNTHESIZED_WIRE_2046 = B[10] & A[3];

assign	SYNTHESIZED_WIRE_2043 = B[10] & A[2];

assign	SYNTHESIZED_WIRE_2040 = B[10] & A[1];

assign	SYNTHESIZED_WIRE_1987 = B[10] & A[0];

assign	SYNTHESIZED_WIRE_1927 = B[11] & A[30];

assign	SYNTHESIZED_WIRE_1930 = ~(A[31] & B[11]);

assign	SYNTHESIZED_WIRE_1924 = B[11] & A[29];


OneBitAdder	b2v_inst138(
	.ci(SYNTHESIZED_WIRE_190),
	.a(SYNTHESIZED_WIRE_191),
	.b(SYNTHESIZED_WIRE_192),
	.co(SYNTHESIZED_WIRE_193),
	.s(SYNTHESIZED_WIRE_94));

assign	SYNTHESIZED_WIRE_1921 = B[11] & A[28];

assign	SYNTHESIZED_WIRE_1918 = B[11] & A[27];

assign	SYNTHESIZED_WIRE_1915 = B[11] & A[26];

assign	SYNTHESIZED_WIRE_1912 = B[11] & A[25];

assign	SYNTHESIZED_WIRE_1909 = B[11] & A[24];

assign	SYNTHESIZED_WIRE_1906 = B[11] & A[23];

assign	SYNTHESIZED_WIRE_1900 = B[11] & A[22];

assign	SYNTHESIZED_WIRE_1897 = B[11] & A[21];

assign	SYNTHESIZED_WIRE_1894 = B[11] & A[20];

assign	SYNTHESIZED_WIRE_1891 = B[11] & A[19];


OneBitAdder	b2v_inst139(
	.ci(SYNTHESIZED_WIRE_193),
	.a(SYNTHESIZED_WIRE_194),
	.b(SYNTHESIZED_WIRE_195),
	.co(SYNTHESIZED_WIRE_196),
	.s(SYNTHESIZED_WIRE_97));

assign	SYNTHESIZED_WIRE_1888 = B[11] & A[18];

assign	SYNTHESIZED_WIRE_1885 = B[11] & A[17];

assign	SYNTHESIZED_WIRE_1984 = B[11] & A[16];

assign	SYNTHESIZED_WIRE_1981 = B[11] & A[15];

assign	SYNTHESIZED_WIRE_1978 = B[11] & A[14];

assign	SYNTHESIZED_WIRE_1975 = B[11] & A[13];

assign	SYNTHESIZED_WIRE_1972 = B[11] & A[12];

assign	SYNTHESIZED_WIRE_1966 = B[11] & A[11];

assign	SYNTHESIZED_WIRE_1963 = B[11] & A[10];

assign	SYNTHESIZED_WIRE_1960 = B[11] & A[9];


OneBitAdder	b2v_inst140(
	.ci(SYNTHESIZED_WIRE_196),
	.a(SYNTHESIZED_WIRE_197),
	.b(SYNTHESIZED_WIRE_198),
	.co(SYNTHESIZED_WIRE_199),
	.s(SYNTHESIZED_WIRE_100));

assign	SYNTHESIZED_WIRE_1957 = B[11] & A[8];

assign	SYNTHESIZED_WIRE_1954 = B[11] & A[7];

assign	SYNTHESIZED_WIRE_1951 = B[11] & A[6];

assign	SYNTHESIZED_WIRE_1948 = B[11] & A[5];

assign	SYNTHESIZED_WIRE_1945 = B[11] & A[4];

assign	SYNTHESIZED_WIRE_1942 = B[11] & A[3];

assign	SYNTHESIZED_WIRE_1939 = B[11] & A[2];

assign	SYNTHESIZED_WIRE_1933 = B[11] & A[1];

assign	SYNTHESIZED_WIRE_1883 = B[11] & A[0];

assign	SYNTHESIZED_WIRE_1823 = B[12] & A[30];


OneBitAdder	b2v_inst141(
	.ci(SYNTHESIZED_WIRE_199),
	.a(SYNTHESIZED_WIRE_200),
	.b(SYNTHESIZED_WIRE_201),
	.co(SYNTHESIZED_WIRE_202),
	.s(SYNTHESIZED_WIRE_103));

assign	SYNTHESIZED_WIRE_1826 = ~(A[31] & B[12]);

assign	SYNTHESIZED_WIRE_1820 = B[12] & A[29];

assign	SYNTHESIZED_WIRE_1817 = B[12] & A[28];

assign	SYNTHESIZED_WIRE_1814 = B[12] & A[27];

assign	SYNTHESIZED_WIRE_1811 = B[12] & A[26];

assign	SYNTHESIZED_WIRE_1808 = B[12] & A[25];

assign	SYNTHESIZED_WIRE_1802 = B[12] & A[24];

assign	SYNTHESIZED_WIRE_1799 = B[12] & A[23];

assign	SYNTHESIZED_WIRE_1796 = B[12] & A[22];

assign	SYNTHESIZED_WIRE_1793 = B[12] & A[21];


OneBitAdder	b2v_inst142(
	.ci(SYNTHESIZED_WIRE_202),
	.a(SYNTHESIZED_WIRE_203),
	.b(SYNTHESIZED_WIRE_204),
	.co(SYNTHESIZED_WIRE_205),
	.s(SYNTHESIZED_WIRE_106));

assign	SYNTHESIZED_WIRE_1790 = B[12] & A[20];

assign	SYNTHESIZED_WIRE_1787 = B[12] & A[19];

assign	SYNTHESIZED_WIRE_1784 = B[12] & A[18];

assign	SYNTHESIZED_WIRE_1781 = B[12] & A[17];

assign	SYNTHESIZED_WIRE_1880 = B[12] & A[16];

assign	SYNTHESIZED_WIRE_1877 = B[12] & A[15];

assign	SYNTHESIZED_WIRE_1874 = B[12] & A[14];

assign	SYNTHESIZED_WIRE_1868 = B[12] & A[13];

assign	SYNTHESIZED_WIRE_1865 = B[12] & A[12];

assign	SYNTHESIZED_WIRE_1862 = B[12] & A[11];


OneBitAdder	b2v_inst143(
	.ci(SYNTHESIZED_WIRE_205),
	.a(SYNTHESIZED_WIRE_206),
	.b(SYNTHESIZED_WIRE_207),
	.co(SYNTHESIZED_WIRE_208),
	.s(SYNTHESIZED_WIRE_109));

assign	SYNTHESIZED_WIRE_1859 = B[12] & A[10];

assign	SYNTHESIZED_WIRE_1856 = B[12] & A[9];

assign	SYNTHESIZED_WIRE_1853 = B[12] & A[8];

assign	SYNTHESIZED_WIRE_1850 = B[12] & A[7];

assign	SYNTHESIZED_WIRE_1847 = B[12] & A[6];

assign	SYNTHESIZED_WIRE_1844 = B[12] & A[5];

assign	SYNTHESIZED_WIRE_1841 = B[12] & A[4];

assign	SYNTHESIZED_WIRE_1835 = B[12] & A[3];

assign	SYNTHESIZED_WIRE_1832 = B[12] & A[2];

assign	SYNTHESIZED_WIRE_1829 = B[12] & A[1];


OneBitAdder	b2v_inst144(
	.ci(SYNTHESIZED_WIRE_208),
	.a(SYNTHESIZED_WIRE_209),
	.b(SYNTHESIZED_WIRE_210),
	.co(SYNTHESIZED_WIRE_115),
	.s(SYNTHESIZED_WIRE_112));

assign	SYNTHESIZED_WIRE_1779 = B[12] & A[0];

assign	SYNTHESIZED_WIRE_1719 = B[13] & A[30];

assign	SYNTHESIZED_WIRE_1722 = ~(A[31] & B[13]);

assign	SYNTHESIZED_WIRE_1716 = B[13] & A[29];

assign	SYNTHESIZED_WIRE_1713 = B[13] & A[28];

assign	SYNTHESIZED_WIRE_1710 = B[13] & A[27];

assign	SYNTHESIZED_WIRE_1704 = B[13] & A[26];

assign	SYNTHESIZED_WIRE_1701 = B[13] & A[25];

assign	SYNTHESIZED_WIRE_1698 = B[13] & A[24];

assign	SYNTHESIZED_WIRE_1695 = B[13] & A[23];


OneBitAdder	b2v_inst145(
	.ci(SYNTHESIZED_WIRE_211),
	.a(SYNTHESIZED_WIRE_212),
	.b(SYNTHESIZED_WIRE_213),
	.co(SYNTHESIZED_WIRE_214),
	.s(SYNTHESIZED_WIRE_2850));

assign	SYNTHESIZED_WIRE_1692 = B[13] & A[22];

assign	SYNTHESIZED_WIRE_1689 = B[13] & A[21];

assign	SYNTHESIZED_WIRE_1686 = B[13] & A[20];

assign	SYNTHESIZED_WIRE_1683 = B[13] & A[19];

assign	SYNTHESIZED_WIRE_1680 = B[13] & A[18];

assign	SYNTHESIZED_WIRE_1677 = B[13] & A[17];

assign	SYNTHESIZED_WIRE_1776 = B[13] & A[16];

assign	SYNTHESIZED_WIRE_1770 = B[13] & A[15];

assign	SYNTHESIZED_WIRE_1767 = B[13] & A[14];

assign	SYNTHESIZED_WIRE_1764 = B[13] & A[13];


OneBitAdder	b2v_inst146(
	.ci(SYNTHESIZED_WIRE_214),
	.a(SYNTHESIZED_WIRE_215),
	.b(SYNTHESIZED_WIRE_216),
	.co(SYNTHESIZED_WIRE_217),
	.s(SYNTHESIZED_WIRE_118));

assign	SYNTHESIZED_WIRE_1761 = B[13] & A[12];

assign	SYNTHESIZED_WIRE_1758 = B[13] & A[11];

assign	SYNTHESIZED_WIRE_1755 = B[13] & A[10];

assign	SYNTHESIZED_WIRE_1752 = B[13] & A[9];

assign	SYNTHESIZED_WIRE_1749 = B[13] & A[8];

assign	SYNTHESIZED_WIRE_1746 = B[13] & A[7];

assign	SYNTHESIZED_WIRE_1743 = B[13] & A[6];

assign	SYNTHESIZED_WIRE_1737 = B[13] & A[5];

assign	SYNTHESIZED_WIRE_1734 = B[13] & A[4];

assign	SYNTHESIZED_WIRE_1731 = B[13] & A[3];


OneBitAdder	b2v_inst147(
	.ci(SYNTHESIZED_WIRE_217),
	.a(SYNTHESIZED_WIRE_218),
	.b(SYNTHESIZED_WIRE_219),
	.co(SYNTHESIZED_WIRE_220),
	.s(SYNTHESIZED_WIRE_121));

assign	SYNTHESIZED_WIRE_1728 = B[13] & A[2];

assign	SYNTHESIZED_WIRE_1725 = B[13] & A[1];

assign	SYNTHESIZED_WIRE_1672 = B[13] & A[0];

assign	SYNTHESIZED_WIRE_1615 = B[14] & A[30];

assign	SYNTHESIZED_WIRE_1618 = ~(A[31] & B[14]);

assign	SYNTHESIZED_WIRE_1612 = B[14] & A[29];

assign	SYNTHESIZED_WIRE_1606 = B[14] & A[28];

assign	SYNTHESIZED_WIRE_1603 = B[14] & A[27];

assign	SYNTHESIZED_WIRE_1600 = B[14] & A[26];

assign	SYNTHESIZED_WIRE_1597 = B[14] & A[25];


OneBitAdder	b2v_inst148(
	.ci(SYNTHESIZED_WIRE_220),
	.a(SYNTHESIZED_WIRE_221),
	.b(SYNTHESIZED_WIRE_222),
	.co(SYNTHESIZED_WIRE_223),
	.s(SYNTHESIZED_WIRE_124));

assign	SYNTHESIZED_WIRE_1594 = B[14] & A[24];

assign	SYNTHESIZED_WIRE_1591 = B[14] & A[23];

assign	SYNTHESIZED_WIRE_1588 = B[14] & A[22];

assign	SYNTHESIZED_WIRE_1585 = B[14] & A[21];

assign	SYNTHESIZED_WIRE_1582 = B[14] & A[20];

assign	SYNTHESIZED_WIRE_1579 = B[14] & A[19];

assign	SYNTHESIZED_WIRE_1573 = B[14] & A[18];

assign	SYNTHESIZED_WIRE_1570 = B[14] & A[17];

assign	SYNTHESIZED_WIRE_1669 = B[14] & A[16];

assign	SYNTHESIZED_WIRE_1666 = B[14] & A[15];


OneBitAdder	b2v_inst149(
	.ci(SYNTHESIZED_WIRE_223),
	.a(SYNTHESIZED_WIRE_224),
	.b(SYNTHESIZED_WIRE_225),
	.co(SYNTHESIZED_WIRE_226),
	.s(SYNTHESIZED_WIRE_127));

assign	SYNTHESIZED_WIRE_1663 = B[14] & A[14];

assign	SYNTHESIZED_WIRE_1660 = B[14] & A[13];

assign	SYNTHESIZED_WIRE_1657 = B[14] & A[12];

assign	SYNTHESIZED_WIRE_1654 = B[14] & A[11];

assign	SYNTHESIZED_WIRE_1651 = B[14] & A[10];

assign	SYNTHESIZED_WIRE_1648 = B[14] & A[9];

assign	SYNTHESIZED_WIRE_1645 = B[14] & A[8];

assign	SYNTHESIZED_WIRE_1639 = B[14] & A[7];

assign	SYNTHESIZED_WIRE_1636 = B[14] & A[6];

assign	SYNTHESIZED_WIRE_1633 = B[14] & A[5];


OneBitAdder	b2v_inst150(
	.ci(SYNTHESIZED_WIRE_226),
	.a(SYNTHESIZED_WIRE_227),
	.b(SYNTHESIZED_WIRE_228),
	.co(SYNTHESIZED_WIRE_229),
	.s(SYNTHESIZED_WIRE_130));

assign	SYNTHESIZED_WIRE_1630 = B[14] & A[4];

assign	SYNTHESIZED_WIRE_1627 = B[14] & A[3];

assign	SYNTHESIZED_WIRE_1624 = B[14] & A[2];

assign	SYNTHESIZED_WIRE_1621 = B[14] & A[1];

assign	SYNTHESIZED_WIRE_1568 = B[14] & A[0];

assign	SYNTHESIZED_WIRE_1508 = B[15] & A[30];

assign	SYNTHESIZED_WIRE_1514 = ~(A[31] & B[15]);

assign	SYNTHESIZED_WIRE_1505 = B[15] & A[29];

assign	SYNTHESIZED_WIRE_1502 = B[15] & A[28];

assign	SYNTHESIZED_WIRE_1499 = B[15] & A[27];


OneBitAdder	b2v_inst151(
	.ci(SYNTHESIZED_WIRE_229),
	.a(SYNTHESIZED_WIRE_230),
	.b(SYNTHESIZED_WIRE_231),
	.co(SYNTHESIZED_WIRE_232),
	.s(SYNTHESIZED_WIRE_133));

assign	SYNTHESIZED_WIRE_1496 = B[15] & A[26];

assign	SYNTHESIZED_WIRE_1493 = B[15] & A[25];

assign	SYNTHESIZED_WIRE_1490 = B[15] & A[24];

assign	SYNTHESIZED_WIRE_1487 = B[15] & A[23];

assign	SYNTHESIZED_WIRE_1484 = B[15] & A[22];

assign	SYNTHESIZED_WIRE_1481 = B[15] & A[21];

assign	SYNTHESIZED_WIRE_1475 = B[15] & A[20];

assign	SYNTHESIZED_WIRE_1472 = B[15] & A[19];

assign	SYNTHESIZED_WIRE_1469 = B[15] & A[18];

assign	SYNTHESIZED_WIRE_1466 = B[15] & A[17];


OneBitAdder	b2v_inst152(
	.ci(SYNTHESIZED_WIRE_232),
	.a(SYNTHESIZED_WIRE_233),
	.b(SYNTHESIZED_WIRE_234),
	.co(SYNTHESIZED_WIRE_235),
	.s(SYNTHESIZED_WIRE_136));

assign	SYNTHESIZED_WIRE_1565 = B[15] & A[16];

assign	SYNTHESIZED_WIRE_1562 = B[15] & A[15];

assign	SYNTHESIZED_WIRE_1559 = B[15] & A[14];

assign	SYNTHESIZED_WIRE_1556 = B[15] & A[13];

assign	SYNTHESIZED_WIRE_1553 = B[15] & A[12];

assign	SYNTHESIZED_WIRE_1550 = B[15] & A[11];

assign	SYNTHESIZED_WIRE_1547 = B[15] & A[10];

assign	SYNTHESIZED_WIRE_1541 = B[15] & A[9];

assign	SYNTHESIZED_WIRE_1538 = B[15] & A[8];

assign	SYNTHESIZED_WIRE_1535 = B[15] & A[7];


OneBitAdder	b2v_inst153(
	.ci(SYNTHESIZED_WIRE_235),
	.a(SYNTHESIZED_WIRE_236),
	.b(SYNTHESIZED_WIRE_237),
	.co(SYNTHESIZED_WIRE_238),
	.s(SYNTHESIZED_WIRE_139));

assign	SYNTHESIZED_WIRE_1532 = B[15] & A[6];

assign	SYNTHESIZED_WIRE_1529 = B[15] & A[5];

assign	SYNTHESIZED_WIRE_1526 = B[15] & A[4];

assign	SYNTHESIZED_WIRE_1523 = B[15] & A[3];

assign	SYNTHESIZED_WIRE_1520 = B[15] & A[2];

assign	SYNTHESIZED_WIRE_1517 = B[15] & A[1];

assign	SYNTHESIZED_WIRE_1464 = B[15] & A[0];

assign	SYNTHESIZED_WIRE_1404 = B[16] & A[30];

assign	SYNTHESIZED_WIRE_1407 = ~(A[31] & B[16]);

assign	SYNTHESIZED_WIRE_1401 = B[16] & A[29];


OneBitAdder	b2v_inst154(
	.ci(SYNTHESIZED_WIRE_238),
	.a(SYNTHESIZED_WIRE_239),
	.b(SYNTHESIZED_WIRE_240),
	.co(SYNTHESIZED_WIRE_241),
	.s(SYNTHESIZED_WIRE_142));

assign	SYNTHESIZED_WIRE_1398 = B[16] & A[28];

assign	SYNTHESIZED_WIRE_1395 = B[16] & A[27];

assign	SYNTHESIZED_WIRE_1392 = B[16] & A[26];

assign	SYNTHESIZED_WIRE_1389 = B[16] & A[25];

assign	SYNTHESIZED_WIRE_1386 = B[16] & A[24];

assign	SYNTHESIZED_WIRE_1383 = B[16] & A[23];

assign	SYNTHESIZED_WIRE_1377 = B[16] & A[22];

assign	SYNTHESIZED_WIRE_1374 = B[16] & A[21];

assign	SYNTHESIZED_WIRE_1371 = B[16] & A[20];

assign	SYNTHESIZED_WIRE_1368 = B[16] & A[19];


OneBitAdder	b2v_inst155(
	.ci(SYNTHESIZED_WIRE_241),
	.a(SYNTHESIZED_WIRE_242),
	.b(SYNTHESIZED_WIRE_243),
	.co(SYNTHESIZED_WIRE_244),
	.s(SYNTHESIZED_WIRE_145));

assign	SYNTHESIZED_WIRE_1365 = B[16] & A[18];

assign	SYNTHESIZED_WIRE_1362 = B[16] & A[17];

assign	SYNTHESIZED_WIRE_1461 = B[16] & A[16];

assign	SYNTHESIZED_WIRE_1458 = B[16] & A[15];

assign	SYNTHESIZED_WIRE_1455 = B[16] & A[14];

assign	SYNTHESIZED_WIRE_1452 = B[16] & A[13];

assign	SYNTHESIZED_WIRE_1449 = B[16] & A[12];

assign	SYNTHESIZED_WIRE_1443 = B[16] & A[11];

assign	SYNTHESIZED_WIRE_1440 = B[16] & A[10];

assign	SYNTHESIZED_WIRE_1437 = B[16] & A[9];


OneBitAdder	b2v_inst156(
	.ci(SYNTHESIZED_WIRE_244),
	.a(SYNTHESIZED_WIRE_245),
	.b(SYNTHESIZED_WIRE_246),
	.co(SYNTHESIZED_WIRE_247),
	.s(SYNTHESIZED_WIRE_148));

assign	SYNTHESIZED_WIRE_1434 = B[16] & A[8];

assign	SYNTHESIZED_WIRE_1431 = B[16] & A[7];

assign	SYNTHESIZED_WIRE_1428 = B[16] & A[6];

assign	SYNTHESIZED_WIRE_1425 = B[16] & A[5];

assign	SYNTHESIZED_WIRE_1422 = B[16] & A[4];

assign	SYNTHESIZED_WIRE_1419 = B[16] & A[3];

assign	SYNTHESIZED_WIRE_1416 = B[16] & A[2];

assign	SYNTHESIZED_WIRE_1410 = B[16] & A[1];

assign	SYNTHESIZED_WIRE_1360 = B[16] & A[0];

assign	SYNTHESIZED_WIRE_1300 = B[17] & A[30];


OneBitAdder	b2v_inst157(
	.ci(SYNTHESIZED_WIRE_247),
	.a(SYNTHESIZED_WIRE_248),
	.b(SYNTHESIZED_WIRE_249),
	.co(SYNTHESIZED_WIRE_250),
	.s(SYNTHESIZED_WIRE_151));

assign	SYNTHESIZED_WIRE_1303 = ~(A[31] & B[17]);

assign	SYNTHESIZED_WIRE_1297 = B[17] & A[29];

assign	SYNTHESIZED_WIRE_1294 = B[17] & A[28];

assign	SYNTHESIZED_WIRE_1291 = B[17] & A[27];

assign	SYNTHESIZED_WIRE_1288 = B[17] & A[26];

assign	SYNTHESIZED_WIRE_1285 = B[17] & A[25];

assign	SYNTHESIZED_WIRE_1279 = B[17] & A[24];

assign	SYNTHESIZED_WIRE_1276 = B[17] & A[23];

assign	SYNTHESIZED_WIRE_1273 = B[17] & A[22];

assign	SYNTHESIZED_WIRE_1270 = B[17] & A[21];


OneBitAdder	b2v_inst158(
	.ci(SYNTHESIZED_WIRE_250),
	.a(SYNTHESIZED_WIRE_251),
	.b(SYNTHESIZED_WIRE_252),
	.co(SYNTHESIZED_WIRE_253),
	.s(SYNTHESIZED_WIRE_154));

assign	SYNTHESIZED_WIRE_1267 = B[17] & A[20];

assign	SYNTHESIZED_WIRE_1264 = B[17] & A[19];

assign	SYNTHESIZED_WIRE_1261 = B[17] & A[18];

assign	SYNTHESIZED_WIRE_1258 = B[17] & A[17];

assign	SYNTHESIZED_WIRE_1357 = B[17] & A[16];

assign	SYNTHESIZED_WIRE_1354 = B[17] & A[15];

assign	SYNTHESIZED_WIRE_1351 = B[17] & A[14];

assign	SYNTHESIZED_WIRE_1345 = B[17] & A[13];

assign	SYNTHESIZED_WIRE_1342 = B[17] & A[12];

assign	SYNTHESIZED_WIRE_1339 = B[17] & A[11];


OneBitAdder	b2v_inst159(
	.ci(SYNTHESIZED_WIRE_253),
	.a(SYNTHESIZED_WIRE_254),
	.b(SYNTHESIZED_WIRE_255),
	.co(SYNTHESIZED_WIRE_256),
	.s(SYNTHESIZED_WIRE_157));

assign	SYNTHESIZED_WIRE_1336 = B[17] & A[10];

assign	SYNTHESIZED_WIRE_1333 = B[17] & A[9];

assign	SYNTHESIZED_WIRE_1330 = B[17] & A[8];

assign	SYNTHESIZED_WIRE_1327 = B[17] & A[7];

assign	SYNTHESIZED_WIRE_1324 = B[17] & A[6];

assign	SYNTHESIZED_WIRE_1321 = B[17] & A[5];

assign	SYNTHESIZED_WIRE_1318 = B[17] & A[4];

assign	SYNTHESIZED_WIRE_1312 = B[17] & A[3];

assign	SYNTHESIZED_WIRE_1309 = B[17] & A[2];

assign	SYNTHESIZED_WIRE_1306 = B[17] & A[1];


OneBitAdder	b2v_inst160(
	.ci(SYNTHESIZED_WIRE_256),
	.a(SYNTHESIZED_WIRE_257),
	.b(SYNTHESIZED_WIRE_258),
	.co(SYNTHESIZED_WIRE_166),
	.s(SYNTHESIZED_WIRE_160));

assign	SYNTHESIZED_WIRE_1256 = B[17] & A[0];

assign	SYNTHESIZED_WIRE_1196 = B[18] & A[30];

assign	SYNTHESIZED_WIRE_1199 = ~(A[31] & B[18]);

assign	SYNTHESIZED_WIRE_1193 = B[18] & A[29];

assign	SYNTHESIZED_WIRE_1190 = B[18] & A[28];

assign	SYNTHESIZED_WIRE_1187 = B[18] & A[27];

assign	SYNTHESIZED_WIRE_1181 = B[18] & A[26];

assign	SYNTHESIZED_WIRE_1178 = B[18] & A[25];

assign	SYNTHESIZED_WIRE_1175 = B[18] & A[24];

assign	SYNTHESIZED_WIRE_1172 = B[18] & A[23];


OneBitAdderHalf	b2v_inst161(
	.A(SYNTHESIZED_WIRE_259),
	.B(SYNTHESIZED_WIRE_260),
	.C(SYNTHESIZED_WIRE_306),
	.S(Z_ALTERA_SYNTHESIZED[27]));

assign	SYNTHESIZED_WIRE_1169 = B[18] & A[22];

assign	SYNTHESIZED_WIRE_1166 = B[18] & A[21];

assign	SYNTHESIZED_WIRE_1163 = B[18] & A[20];

assign	SYNTHESIZED_WIRE_1160 = B[18] & A[19];

assign	SYNTHESIZED_WIRE_1157 = B[18] & A[18];

assign	SYNTHESIZED_WIRE_1154 = B[18] & A[17];

assign	SYNTHESIZED_WIRE_1253 = B[18] & A[16];

assign	SYNTHESIZED_WIRE_1247 = B[18] & A[15];

assign	SYNTHESIZED_WIRE_1244 = B[18] & A[14];

assign	SYNTHESIZED_WIRE_1241 = B[18] & A[13];


OneBitAdder	b2v_inst162(
	.ci(SYNTHESIZED_WIRE_261),
	.a(SYNTHESIZED_WIRE_262),
	.b(SYNTHESIZED_WIRE_263),
	.co(SYNTHESIZED_WIRE_264),
	.s(SYNTHESIZED_WIRE_258));

assign	SYNTHESIZED_WIRE_1238 = B[18] & A[12];

assign	SYNTHESIZED_WIRE_1235 = B[18] & A[11];

assign	SYNTHESIZED_WIRE_1232 = B[18] & A[10];

assign	SYNTHESIZED_WIRE_1229 = B[18] & A[9];

assign	SYNTHESIZED_WIRE_1226 = B[18] & A[8];

assign	SYNTHESIZED_WIRE_1223 = B[18] & A[7];

assign	SYNTHESIZED_WIRE_1220 = B[18] & A[6];

assign	SYNTHESIZED_WIRE_1214 = B[18] & A[5];

assign	SYNTHESIZED_WIRE_1211 = B[18] & A[4];

assign	SYNTHESIZED_WIRE_1208 = B[18] & A[3];


OneBitAdder	b2v_inst163(
	.ci(SYNTHESIZED_WIRE_264),
	.a(SYNTHESIZED_WIRE_265),
	.b(SYNTHESIZED_WIRE_266),
	.co(SYNTHESIZED_WIRE_267),
	.s(SYNTHESIZED_WIRE_168));

assign	SYNTHESIZED_WIRE_1205 = B[18] & A[2];

assign	SYNTHESIZED_WIRE_1202 = B[18] & A[1];

assign	SYNTHESIZED_WIRE_1149 = B[18] & A[0];

assign	SYNTHESIZED_WIRE_1092 = B[19] & A[30];

assign	SYNTHESIZED_WIRE_1095 = ~(A[31] & B[19]);

assign	SYNTHESIZED_WIRE_1089 = B[19] & A[29];

assign	SYNTHESIZED_WIRE_1083 = B[19] & A[28];

assign	SYNTHESIZED_WIRE_1080 = B[19] & A[27];

assign	SYNTHESIZED_WIRE_1077 = B[19] & A[26];

assign	SYNTHESIZED_WIRE_1074 = B[19] & A[25];


OneBitAdder	b2v_inst164(
	.ci(SYNTHESIZED_WIRE_267),
	.a(SYNTHESIZED_WIRE_268),
	.b(SYNTHESIZED_WIRE_269),
	.co(SYNTHESIZED_WIRE_270),
	.s(SYNTHESIZED_WIRE_171));

assign	SYNTHESIZED_WIRE_1071 = B[19] & A[24];

assign	SYNTHESIZED_WIRE_1068 = B[19] & A[23];

assign	SYNTHESIZED_WIRE_1065 = B[19] & A[22];

assign	SYNTHESIZED_WIRE_1062 = B[19] & A[21];

assign	SYNTHESIZED_WIRE_1059 = B[19] & A[20];

assign	SYNTHESIZED_WIRE_1056 = B[19] & A[19];

assign	SYNTHESIZED_WIRE_1050 = B[19] & A[18];

assign	SYNTHESIZED_WIRE_1047 = B[19] & A[17];

assign	SYNTHESIZED_WIRE_1146 = B[19] & A[16];

assign	SYNTHESIZED_WIRE_1143 = B[19] & A[15];


OneBitAdder	b2v_inst165(
	.ci(SYNTHESIZED_WIRE_270),
	.a(SYNTHESIZED_WIRE_271),
	.b(SYNTHESIZED_WIRE_272),
	.co(SYNTHESIZED_WIRE_273),
	.s(SYNTHESIZED_WIRE_174));

assign	SYNTHESIZED_WIRE_1140 = B[19] & A[14];

assign	SYNTHESIZED_WIRE_1137 = B[19] & A[13];

assign	SYNTHESIZED_WIRE_1134 = B[19] & A[12];

assign	SYNTHESIZED_WIRE_1131 = B[19] & A[11];

assign	SYNTHESIZED_WIRE_1128 = B[19] & A[10];

assign	SYNTHESIZED_WIRE_1125 = B[19] & A[9];

assign	SYNTHESIZED_WIRE_1122 = B[19] & A[8];

assign	SYNTHESIZED_WIRE_1116 = B[19] & A[7];

assign	SYNTHESIZED_WIRE_1113 = B[19] & A[6];

assign	SYNTHESIZED_WIRE_1110 = B[19] & A[5];


OneBitAdder	b2v_inst166(
	.ci(SYNTHESIZED_WIRE_273),
	.a(SYNTHESIZED_WIRE_274),
	.b(SYNTHESIZED_WIRE_275),
	.co(SYNTHESIZED_WIRE_276),
	.s(SYNTHESIZED_WIRE_177));

assign	SYNTHESIZED_WIRE_1107 = B[19] & A[4];

assign	SYNTHESIZED_WIRE_1104 = B[19] & A[3];

assign	SYNTHESIZED_WIRE_1101 = B[19] & A[2];

assign	SYNTHESIZED_WIRE_1098 = B[19] & A[1];

assign	SYNTHESIZED_WIRE_1045 = B[19] & A[0];

assign	SYNTHESIZED_WIRE_985 = B[20] & A[30];

assign	SYNTHESIZED_WIRE_991 = ~(A[31] & B[20]);

assign	SYNTHESIZED_WIRE_982 = B[20] & A[29];

assign	SYNTHESIZED_WIRE_979 = B[20] & A[28];

assign	SYNTHESIZED_WIRE_976 = B[20] & A[27];


OneBitAdder	b2v_inst167(
	.ci(SYNTHESIZED_WIRE_276),
	.a(SYNTHESIZED_WIRE_277),
	.b(SYNTHESIZED_WIRE_278),
	.co(SYNTHESIZED_WIRE_279),
	.s(SYNTHESIZED_WIRE_180));

assign	SYNTHESIZED_WIRE_973 = B[20] & A[26];

assign	SYNTHESIZED_WIRE_970 = B[20] & A[25];

assign	SYNTHESIZED_WIRE_967 = B[20] & A[24];

assign	SYNTHESIZED_WIRE_964 = B[20] & A[23];

assign	SYNTHESIZED_WIRE_961 = B[20] & A[22];

assign	SYNTHESIZED_WIRE_958 = B[20] & A[21];

assign	SYNTHESIZED_WIRE_952 = B[20] & A[20];

assign	SYNTHESIZED_WIRE_949 = B[20] & A[19];

assign	SYNTHESIZED_WIRE_946 = B[20] & A[18];

assign	SYNTHESIZED_WIRE_943 = B[20] & A[17];


OneBitAdder	b2v_inst168(
	.ci(SYNTHESIZED_WIRE_279),
	.a(SYNTHESIZED_WIRE_280),
	.b(SYNTHESIZED_WIRE_281),
	.co(SYNTHESIZED_WIRE_282),
	.s(SYNTHESIZED_WIRE_183));

assign	SYNTHESIZED_WIRE_1042 = B[20] & A[16];

assign	SYNTHESIZED_WIRE_1039 = B[20] & A[15];

assign	SYNTHESIZED_WIRE_1036 = B[20] & A[14];

assign	SYNTHESIZED_WIRE_1033 = B[20] & A[13];

assign	SYNTHESIZED_WIRE_1030 = B[20] & A[12];

assign	SYNTHESIZED_WIRE_1027 = B[20] & A[11];

assign	SYNTHESIZED_WIRE_1024 = B[20] & A[10];

assign	SYNTHESIZED_WIRE_1018 = B[20] & A[9];

assign	SYNTHESIZED_WIRE_1015 = B[20] & A[8];

assign	SYNTHESIZED_WIRE_1012 = B[20] & A[7];


OneBitAdder	b2v_inst169(
	.ci(SYNTHESIZED_WIRE_282),
	.a(SYNTHESIZED_WIRE_283),
	.b(SYNTHESIZED_WIRE_284),
	.co(SYNTHESIZED_WIRE_285),
	.s(SYNTHESIZED_WIRE_186));

assign	SYNTHESIZED_WIRE_1009 = B[20] & A[6];

assign	SYNTHESIZED_WIRE_1006 = B[20] & A[5];

assign	SYNTHESIZED_WIRE_1003 = B[20] & A[4];

assign	SYNTHESIZED_WIRE_1000 = B[20] & A[3];

assign	SYNTHESIZED_WIRE_997 = B[20] & A[2];

assign	SYNTHESIZED_WIRE_994 = B[20] & A[1];

assign	SYNTHESIZED_WIRE_941 = B[20] & A[0];

assign	SYNTHESIZED_WIRE_881 = B[21] & A[30];

assign	SYNTHESIZED_WIRE_884 = ~(A[31] & B[21]);

assign	SYNTHESIZED_WIRE_878 = B[21] & A[29];


OneBitAdder	b2v_inst170(
	.ci(SYNTHESIZED_WIRE_285),
	.a(SYNTHESIZED_WIRE_286),
	.b(SYNTHESIZED_WIRE_287),
	.co(SYNTHESIZED_WIRE_288),
	.s(SYNTHESIZED_WIRE_189));

assign	SYNTHESIZED_WIRE_875 = B[21] & A[28];

assign	SYNTHESIZED_WIRE_872 = B[21] & A[27];

assign	SYNTHESIZED_WIRE_869 = B[21] & A[26];

assign	SYNTHESIZED_WIRE_866 = B[21] & A[25];

assign	SYNTHESIZED_WIRE_863 = B[21] & A[24];

assign	SYNTHESIZED_WIRE_860 = B[21] & A[23];

assign	SYNTHESIZED_WIRE_854 = B[21] & A[22];

assign	SYNTHESIZED_WIRE_851 = B[21] & A[21];

assign	SYNTHESIZED_WIRE_848 = B[21] & A[20];

assign	SYNTHESIZED_WIRE_845 = B[21] & A[19];


OneBitAdder	b2v_inst171(
	.ci(SYNTHESIZED_WIRE_288),
	.a(SYNTHESIZED_WIRE_289),
	.b(SYNTHESIZED_WIRE_290),
	.co(SYNTHESIZED_WIRE_291),
	.s(SYNTHESIZED_WIRE_192));

assign	SYNTHESIZED_WIRE_842 = B[21] & A[18];

assign	SYNTHESIZED_WIRE_839 = B[21] & A[17];

assign	SYNTHESIZED_WIRE_938 = B[21] & A[16];

assign	SYNTHESIZED_WIRE_935 = B[21] & A[15];

assign	SYNTHESIZED_WIRE_932 = B[21] & A[14];

assign	SYNTHESIZED_WIRE_929 = B[21] & A[13];

assign	SYNTHESIZED_WIRE_926 = B[21] & A[12];

assign	SYNTHESIZED_WIRE_920 = B[21] & A[11];

assign	SYNTHESIZED_WIRE_917 = B[21] & A[10];

assign	SYNTHESIZED_WIRE_914 = B[21] & A[9];


OneBitAdder	b2v_inst172(
	.ci(SYNTHESIZED_WIRE_291),
	.a(SYNTHESIZED_WIRE_292),
	.b(SYNTHESIZED_WIRE_293),
	.co(SYNTHESIZED_WIRE_294),
	.s(SYNTHESIZED_WIRE_195));

assign	SYNTHESIZED_WIRE_911 = B[21] & A[8];

assign	SYNTHESIZED_WIRE_908 = B[21] & A[7];

assign	SYNTHESIZED_WIRE_905 = B[21] & A[6];

assign	SYNTHESIZED_WIRE_902 = B[21] & A[5];

assign	SYNTHESIZED_WIRE_899 = B[21] & A[4];

assign	SYNTHESIZED_WIRE_896 = B[21] & A[3];

assign	SYNTHESIZED_WIRE_893 = B[21] & A[2];

assign	SYNTHESIZED_WIRE_887 = B[21] & A[1];

assign	SYNTHESIZED_WIRE_837 = B[21] & A[0];

assign	SYNTHESIZED_WIRE_780 = B[22] & A[30];


OneBitAdder	b2v_inst173(
	.ci(SYNTHESIZED_WIRE_294),
	.a(SYNTHESIZED_WIRE_295),
	.b(SYNTHESIZED_WIRE_296),
	.co(SYNTHESIZED_WIRE_297),
	.s(SYNTHESIZED_WIRE_198));

assign	SYNTHESIZED_WIRE_783 = ~(A[31] & B[22]);

assign	SYNTHESIZED_WIRE_777 = B[22] & A[29];

assign	SYNTHESIZED_WIRE_774 = B[22] & A[28];

assign	SYNTHESIZED_WIRE_771 = B[22] & A[27];

assign	SYNTHESIZED_WIRE_768 = B[22] & A[26];

assign	SYNTHESIZED_WIRE_765 = B[22] & A[25];

assign	SYNTHESIZED_WIRE_762 = B[22] & A[24];

assign	SYNTHESIZED_WIRE_759 = B[22] & A[23];

assign	SYNTHESIZED_WIRE_756 = B[22] & A[22];

assign	SYNTHESIZED_WIRE_753 = B[22] & A[21];


OneBitAdder	b2v_inst174(
	.ci(SYNTHESIZED_WIRE_297),
	.a(SYNTHESIZED_WIRE_298),
	.b(SYNTHESIZED_WIRE_299),
	.co(SYNTHESIZED_WIRE_300),
	.s(SYNTHESIZED_WIRE_201));

assign	SYNTHESIZED_WIRE_750 = B[22] & A[20];

assign	SYNTHESIZED_WIRE_747 = B[22] & A[19];

assign	SYNTHESIZED_WIRE_744 = B[22] & A[18];

assign	SYNTHESIZED_WIRE_741 = B[22] & A[17];

assign	SYNTHESIZED_WIRE_834 = B[22] & A[16];

assign	SYNTHESIZED_WIRE_831 = B[22] & A[15];

assign	SYNTHESIZED_WIRE_828 = B[22] & A[14];

assign	SYNTHESIZED_WIRE_822 = B[22] & A[13];

assign	SYNTHESIZED_WIRE_819 = B[22] & A[12];

assign	SYNTHESIZED_WIRE_816 = B[22] & A[11];


OneBitAdder	b2v_inst175(
	.ci(SYNTHESIZED_WIRE_300),
	.a(SYNTHESIZED_WIRE_301),
	.b(SYNTHESIZED_WIRE_302),
	.co(SYNTHESIZED_WIRE_303),
	.s(SYNTHESIZED_WIRE_204));

assign	SYNTHESIZED_WIRE_813 = B[22] & A[10];

assign	SYNTHESIZED_WIRE_810 = B[22] & A[9];

assign	SYNTHESIZED_WIRE_807 = B[22] & A[8];

assign	SYNTHESIZED_WIRE_804 = B[22] & A[7];

assign	SYNTHESIZED_WIRE_801 = B[22] & A[6];

assign	SYNTHESIZED_WIRE_798 = B[22] & A[5];

assign	SYNTHESIZED_WIRE_795 = B[22] & A[4];

assign	SYNTHESIZED_WIRE_792 = B[22] & A[3];

assign	SYNTHESIZED_WIRE_789 = B[22] & A[2];

assign	SYNTHESIZED_WIRE_786 = B[22] & A[1];


OneBitAdder	b2v_inst176(
	.ci(SYNTHESIZED_WIRE_303),
	.a(SYNTHESIZED_WIRE_304),
	.b(SYNTHESIZED_WIRE_305),
	.co(SYNTHESIZED_WIRE_210),
	.s(SYNTHESIZED_WIRE_207));

assign	SYNTHESIZED_WIRE_739 = B[22] & A[0];

assign	SYNTHESIZED_WIRE_685 = B[23] & A[30];

assign	SYNTHESIZED_WIRE_688 = ~(A[31] & B[23]);

assign	SYNTHESIZED_WIRE_682 = B[23] & A[29];

assign	SYNTHESIZED_WIRE_679 = B[23] & A[28];

assign	SYNTHESIZED_WIRE_676 = B[23] & A[27];

assign	SYNTHESIZED_WIRE_671 = B[23] & A[26];

assign	SYNTHESIZED_WIRE_668 = B[23] & A[25];

assign	SYNTHESIZED_WIRE_665 = B[23] & A[24];

assign	SYNTHESIZED_WIRE_662 = B[23] & A[23];


OneBitAdder	b2v_inst177(
	.ci(SYNTHESIZED_WIRE_306),
	.a(SYNTHESIZED_WIRE_307),
	.b(SYNTHESIZED_WIRE_308),
	.co(SYNTHESIZED_WIRE_309),
	.s(SYNTHESIZED_WIRE_164));

assign	SYNTHESIZED_WIRE_659 = B[23] & A[22];

assign	SYNTHESIZED_WIRE_656 = B[23] & A[21];

assign	SYNTHESIZED_WIRE_653 = B[23] & A[20];

assign	SYNTHESIZED_WIRE_650 = B[23] & A[19];

assign	SYNTHESIZED_WIRE_647 = B[23] & A[18];

assign	SYNTHESIZED_WIRE_644 = B[23] & A[17];

assign	SYNTHESIZED_WIRE_736 = B[23] & A[16];

assign	SYNTHESIZED_WIRE_733 = B[23] & A[15];

assign	SYNTHESIZED_WIRE_730 = B[23] & A[14];

assign	SYNTHESIZED_WIRE_727 = B[23] & A[13];


OneBitAdder	b2v_inst178(
	.ci(SYNTHESIZED_WIRE_309),
	.a(SYNTHESIZED_WIRE_310),
	.b(SYNTHESIZED_WIRE_311),
	.co(SYNTHESIZED_WIRE_312),
	.s(SYNTHESIZED_WIRE_213));

assign	SYNTHESIZED_WIRE_724 = B[23] & A[12];

assign	SYNTHESIZED_WIRE_721 = B[23] & A[11];

assign	SYNTHESIZED_WIRE_718 = B[23] & A[10];

assign	SYNTHESIZED_WIRE_715 = B[23] & A[9];

assign	SYNTHESIZED_WIRE_712 = B[23] & A[8];

assign	SYNTHESIZED_WIRE_709 = B[23] & A[7];

assign	SYNTHESIZED_WIRE_706 = B[23] & A[6];

assign	SYNTHESIZED_WIRE_703 = B[23] & A[5];

assign	SYNTHESIZED_WIRE_700 = B[23] & A[4];

assign	SYNTHESIZED_WIRE_697 = B[23] & A[3];


OneBitAdder	b2v_inst179(
	.ci(SYNTHESIZED_WIRE_312),
	.a(SYNTHESIZED_WIRE_313),
	.b(SYNTHESIZED_WIRE_314),
	.co(SYNTHESIZED_WIRE_315),
	.s(SYNTHESIZED_WIRE_216));

assign	SYNTHESIZED_WIRE_694 = B[23] & A[2];

assign	SYNTHESIZED_WIRE_691 = B[23] & A[1];

assign	SYNTHESIZED_WIRE_642 = B[23] & A[0];

assign	SYNTHESIZED_WIRE_588 = B[24] & A[30];

assign	SYNTHESIZED_WIRE_591 = ~(A[31] & B[24]);

assign	SYNTHESIZED_WIRE_585 = B[24] & A[29];

assign	SYNTHESIZED_WIRE_582 = B[24] & A[28];

assign	SYNTHESIZED_WIRE_579 = B[24] & A[27];

assign	SYNTHESIZED_WIRE_576 = B[24] & A[26];

assign	SYNTHESIZED_WIRE_573 = B[24] & A[25];


OneBitAdder	b2v_inst180(
	.ci(SYNTHESIZED_WIRE_315),
	.a(SYNTHESIZED_WIRE_316),
	.b(SYNTHESIZED_WIRE_317),
	.co(SYNTHESIZED_WIRE_318),
	.s(SYNTHESIZED_WIRE_219));

assign	SYNTHESIZED_WIRE_570 = B[24] & A[24];

assign	SYNTHESIZED_WIRE_567 = B[24] & A[23];

assign	SYNTHESIZED_WIRE_564 = B[24] & A[22];

assign	SYNTHESIZED_WIRE_561 = B[24] & A[21];

assign	SYNTHESIZED_WIRE_558 = B[24] & A[20];

assign	SYNTHESIZED_WIRE_555 = B[24] & A[19];

assign	SYNTHESIZED_WIRE_552 = B[24] & A[18];

assign	SYNTHESIZED_WIRE_549 = B[24] & A[17];

assign	SYNTHESIZED_WIRE_639 = B[24] & A[16];

assign	SYNTHESIZED_WIRE_636 = B[24] & A[15];


OneBitAdder	b2v_inst181(
	.ci(SYNTHESIZED_WIRE_318),
	.a(SYNTHESIZED_WIRE_319),
	.b(SYNTHESIZED_WIRE_320),
	.co(SYNTHESIZED_WIRE_321),
	.s(SYNTHESIZED_WIRE_222));

assign	SYNTHESIZED_WIRE_633 = B[24] & A[14];

assign	SYNTHESIZED_WIRE_630 = B[24] & A[13];

assign	SYNTHESIZED_WIRE_627 = B[24] & A[12];

assign	SYNTHESIZED_WIRE_624 = B[24] & A[11];

assign	SYNTHESIZED_WIRE_621 = B[24] & A[10];

assign	SYNTHESIZED_WIRE_618 = B[24] & A[9];

assign	SYNTHESIZED_WIRE_615 = B[24] & A[8];

assign	SYNTHESIZED_WIRE_612 = B[24] & A[7];

assign	SYNTHESIZED_WIRE_609 = B[24] & A[6];

assign	SYNTHESIZED_WIRE_606 = B[24] & A[5];


OneBitAdder	b2v_inst182(
	.ci(SYNTHESIZED_WIRE_321),
	.a(SYNTHESIZED_WIRE_322),
	.b(SYNTHESIZED_WIRE_323),
	.co(SYNTHESIZED_WIRE_324),
	.s(SYNTHESIZED_WIRE_225));

assign	SYNTHESIZED_WIRE_603 = B[24] & A[4];

assign	SYNTHESIZED_WIRE_600 = B[24] & A[3];

assign	SYNTHESIZED_WIRE_597 = B[24] & A[2];

assign	SYNTHESIZED_WIRE_594 = B[24] & A[1];

assign	SYNTHESIZED_WIRE_547 = B[24] & A[0];

assign	SYNTHESIZED_WIRE_493 = B[25] & A[30];

assign	SYNTHESIZED_WIRE_496 = ~(A[31] & B[25]);

assign	SYNTHESIZED_WIRE_490 = B[25] & A[29];

assign	SYNTHESIZED_WIRE_487 = B[25] & A[28];

assign	SYNTHESIZED_WIRE_484 = B[25] & A[27];


OneBitAdder	b2v_inst183(
	.ci(SYNTHESIZED_WIRE_324),
	.a(SYNTHESIZED_WIRE_325),
	.b(SYNTHESIZED_WIRE_326),
	.co(SYNTHESIZED_WIRE_327),
	.s(SYNTHESIZED_WIRE_228));

assign	SYNTHESIZED_WIRE_481 = B[25] & A[26];

assign	SYNTHESIZED_WIRE_478 = B[25] & A[25];

assign	SYNTHESIZED_WIRE_475 = B[25] & A[24];

assign	SYNTHESIZED_WIRE_472 = B[25] & A[23];

assign	SYNTHESIZED_WIRE_469 = B[25] & A[22];

assign	SYNTHESIZED_WIRE_466 = B[25] & A[21];

assign	SYNTHESIZED_WIRE_463 = B[25] & A[20];

assign	SYNTHESIZED_WIRE_460 = B[25] & A[19];

assign	SYNTHESIZED_WIRE_457 = B[25] & A[18];

assign	SYNTHESIZED_WIRE_454 = B[25] & A[17];


OneBitAdder	b2v_inst184(
	.ci(SYNTHESIZED_WIRE_327),
	.a(SYNTHESIZED_WIRE_328),
	.b(SYNTHESIZED_WIRE_329),
	.co(SYNTHESIZED_WIRE_330),
	.s(SYNTHESIZED_WIRE_231));

assign	SYNTHESIZED_WIRE_544 = B[25] & A[16];

assign	SYNTHESIZED_WIRE_541 = B[25] & A[15];

assign	SYNTHESIZED_WIRE_538 = B[25] & A[14];

assign	SYNTHESIZED_WIRE_535 = B[25] & A[13];

assign	SYNTHESIZED_WIRE_532 = B[25] & A[12];

assign	SYNTHESIZED_WIRE_529 = B[25] & A[11];

assign	SYNTHESIZED_WIRE_526 = B[25] & A[10];

assign	SYNTHESIZED_WIRE_523 = B[25] & A[9];

assign	SYNTHESIZED_WIRE_520 = B[25] & A[8];

assign	SYNTHESIZED_WIRE_517 = B[25] & A[7];


OneBitAdder	b2v_inst185(
	.ci(SYNTHESIZED_WIRE_330),
	.a(SYNTHESIZED_WIRE_331),
	.b(SYNTHESIZED_WIRE_332),
	.co(SYNTHESIZED_WIRE_333),
	.s(SYNTHESIZED_WIRE_234));

assign	SYNTHESIZED_WIRE_514 = B[25] & A[6];

assign	SYNTHESIZED_WIRE_511 = B[25] & A[5];

assign	SYNTHESIZED_WIRE_508 = B[25] & A[4];

assign	SYNTHESIZED_WIRE_505 = B[25] & A[3];

assign	SYNTHESIZED_WIRE_502 = B[25] & A[2];

assign	SYNTHESIZED_WIRE_499 = B[25] & A[1];

assign	SYNTHESIZED_WIRE_452 = B[25] & A[0];

assign	SYNTHESIZED_WIRE_1282 = B[31] & A[31];


OneBitAdder	b2v_inst186(
	.ci(SYNTHESIZED_WIRE_333),
	.a(SYNTHESIZED_WIRE_334),
	.b(SYNTHESIZED_WIRE_335),
	.co(SYNTHESIZED_WIRE_336),
	.s(SYNTHESIZED_WIRE_237));


OneBitAdder	b2v_inst187(
	.ci(SYNTHESIZED_WIRE_336),
	.a(SYNTHESIZED_WIRE_337),
	.b(SYNTHESIZED_WIRE_338),
	.co(SYNTHESIZED_WIRE_339),
	.s(SYNTHESIZED_WIRE_240));


OneBitAdder	b2v_inst188(
	.ci(SYNTHESIZED_WIRE_339),
	.a(SYNTHESIZED_WIRE_340),
	.b(SYNTHESIZED_WIRE_341),
	.co(SYNTHESIZED_WIRE_342),
	.s(SYNTHESIZED_WIRE_243));

assign	SYNTHESIZED_WIRE_1 = ~(A[0] & B[31]);



OneBitAdder	b2v_inst189(
	.ci(SYNTHESIZED_WIRE_342),
	.a(SYNTHESIZED_WIRE_343),
	.b(SYNTHESIZED_WIRE_344),
	.co(SYNTHESIZED_WIRE_345),
	.s(SYNTHESIZED_WIRE_246));

assign	SYNTHESIZED_WIRE_398 = B[26] & A[30];

assign	SYNTHESIZED_WIRE_401 = ~(A[31] & B[26]);

assign	SYNTHESIZED_WIRE_395 = B[26] & A[29];

assign	SYNTHESIZED_WIRE_392 = B[26] & A[28];

assign	SYNTHESIZED_WIRE_389 = B[26] & A[27];

assign	SYNTHESIZED_WIRE_386 = B[26] & A[26];

assign	SYNTHESIZED_WIRE_383 = B[26] & A[25];

assign	SYNTHESIZED_WIRE_380 = B[26] & A[24];

assign	SYNTHESIZED_WIRE_377 = B[26] & A[23];

assign	SYNTHESIZED_WIRE_372 = B[26] & A[22];


OneBitAdder	b2v_inst190(
	.ci(SYNTHESIZED_WIRE_345),
	.a(SYNTHESIZED_WIRE_346),
	.b(SYNTHESIZED_WIRE_347),
	.co(SYNTHESIZED_WIRE_348),
	.s(SYNTHESIZED_WIRE_249));

assign	SYNTHESIZED_WIRE_369 = B[26] & A[21];

assign	SYNTHESIZED_WIRE_366 = B[26] & A[20];

assign	SYNTHESIZED_WIRE_363 = B[26] & A[19];

assign	SYNTHESIZED_WIRE_360 = B[26] & A[18];

assign	SYNTHESIZED_WIRE_357 = B[26] & A[17];

assign	SYNTHESIZED_WIRE_449 = B[26] & A[16];

assign	SYNTHESIZED_WIRE_446 = B[26] & A[15];

assign	SYNTHESIZED_WIRE_443 = B[26] & A[14];

assign	SYNTHESIZED_WIRE_440 = B[26] & A[13];

assign	SYNTHESIZED_WIRE_437 = B[26] & A[12];


OneBitAdder	b2v_inst191(
	.ci(SYNTHESIZED_WIRE_348),
	.a(SYNTHESIZED_WIRE_349),
	.b(SYNTHESIZED_WIRE_350),
	.co(SYNTHESIZED_WIRE_351),
	.s(SYNTHESIZED_WIRE_252));

assign	SYNTHESIZED_WIRE_434 = B[26] & A[11];

assign	SYNTHESIZED_WIRE_431 = B[26] & A[10];

assign	SYNTHESIZED_WIRE_428 = B[26] & A[9];

assign	SYNTHESIZED_WIRE_425 = B[26] & A[8];

assign	SYNTHESIZED_WIRE_422 = B[26] & A[7];

assign	SYNTHESIZED_WIRE_419 = B[26] & A[6];

assign	SYNTHESIZED_WIRE_416 = B[26] & A[5];

assign	SYNTHESIZED_WIRE_413 = B[26] & A[4];

assign	SYNTHESIZED_WIRE_410 = B[26] & A[3];

assign	SYNTHESIZED_WIRE_407 = B[26] & A[2];


OneBitAdder	b2v_inst192(
	.ci(SYNTHESIZED_WIRE_351),
	.a(SYNTHESIZED_WIRE_352),
	.b(SYNTHESIZED_WIRE_353),
	.co(SYNTHESIZED_WIRE_261),
	.s(SYNTHESIZED_WIRE_255));

assign	SYNTHESIZED_WIRE_404 = B[26] & A[1];

assign	SYNTHESIZED_WIRE_355 = B[26] & A[0];

assign	SYNTHESIZED_WIRE_301 = B[27] & A[30];

assign	SYNTHESIZED_WIRE_304 = ~(A[31] & B[27]);

assign	SYNTHESIZED_WIRE_298 = B[27] & A[29];

assign	SYNTHESIZED_WIRE_295 = B[27] & A[28];

assign	SYNTHESIZED_WIRE_292 = B[27] & A[27];

assign	SYNTHESIZED_WIRE_289 = B[27] & A[26];

assign	SYNTHESIZED_WIRE_286 = B[27] & A[25];

assign	SYNTHESIZED_WIRE_283 = B[27] & A[24];


OneBitAdderHalf	b2v_inst193(
	.A(SYNTHESIZED_WIRE_354),
	.B(SYNTHESIZED_WIRE_355),
	.C(SYNTHESIZED_WIRE_403),
	.S(Z_ALTERA_SYNTHESIZED[26]));

assign	SYNTHESIZED_WIRE_280 = B[27] & A[23];

assign	SYNTHESIZED_WIRE_277 = B[27] & A[22];

assign	SYNTHESIZED_WIRE_274 = B[27] & A[21];

assign	SYNTHESIZED_WIRE_271 = B[27] & A[20];

assign	SYNTHESIZED_WIRE_268 = B[27] & A[19];

assign	SYNTHESIZED_WIRE_265 = B[27] & A[18];

assign	SYNTHESIZED_WIRE_262 = B[27] & A[17];

assign	SYNTHESIZED_WIRE_352 = B[27] & A[16];

assign	SYNTHESIZED_WIRE_349 = B[27] & A[15];

assign	SYNTHESIZED_WIRE_346 = B[27] & A[14];


OneBitAdder	b2v_inst194(
	.ci(SYNTHESIZED_WIRE_356),
	.a(SYNTHESIZED_WIRE_357),
	.b(SYNTHESIZED_WIRE_358),
	.co(SYNTHESIZED_WIRE_359),
	.s(SYNTHESIZED_WIRE_353));

assign	SYNTHESIZED_WIRE_343 = B[27] & A[13];

assign	SYNTHESIZED_WIRE_340 = B[27] & A[12];

assign	SYNTHESIZED_WIRE_337 = B[27] & A[11];

assign	SYNTHESIZED_WIRE_334 = B[27] & A[10];

assign	SYNTHESIZED_WIRE_331 = B[27] & A[9];

assign	SYNTHESIZED_WIRE_328 = B[27] & A[8];

assign	SYNTHESIZED_WIRE_325 = B[27] & A[7];

assign	SYNTHESIZED_WIRE_322 = B[27] & A[6];

assign	SYNTHESIZED_WIRE_319 = B[27] & A[5];

assign	SYNTHESIZED_WIRE_316 = B[27] & A[4];


OneBitAdder	b2v_inst195(
	.ci(SYNTHESIZED_WIRE_359),
	.a(SYNTHESIZED_WIRE_360),
	.b(SYNTHESIZED_WIRE_361),
	.co(SYNTHESIZED_WIRE_362),
	.s(SYNTHESIZED_WIRE_263));

assign	SYNTHESIZED_WIRE_313 = B[27] & A[3];

assign	SYNTHESIZED_WIRE_310 = B[27] & A[2];

assign	SYNTHESIZED_WIRE_307 = B[27] & A[1];

assign	SYNTHESIZED_WIRE_260 = B[27] & A[0];

assign	SYNTHESIZED_WIRE_206 = B[28] & A[30];

assign	SYNTHESIZED_WIRE_209 = ~(A[31] & B[28]);

assign	SYNTHESIZED_WIRE_203 = B[28] & A[29];

assign	SYNTHESIZED_WIRE_200 = B[28] & A[28];

assign	SYNTHESIZED_WIRE_197 = B[28] & A[27];

assign	SYNTHESIZED_WIRE_194 = B[28] & A[26];


OneBitAdder	b2v_inst196(
	.ci(SYNTHESIZED_WIRE_362),
	.a(SYNTHESIZED_WIRE_363),
	.b(SYNTHESIZED_WIRE_364),
	.co(SYNTHESIZED_WIRE_365),
	.s(SYNTHESIZED_WIRE_266));

assign	SYNTHESIZED_WIRE_191 = B[28] & A[25];

assign	SYNTHESIZED_WIRE_188 = B[28] & A[24];

assign	SYNTHESIZED_WIRE_185 = B[28] & A[23];

assign	SYNTHESIZED_WIRE_182 = B[28] & A[22];

assign	SYNTHESIZED_WIRE_179 = B[28] & A[21];

assign	SYNTHESIZED_WIRE_176 = B[28] & A[20];

assign	SYNTHESIZED_WIRE_173 = B[28] & A[19];

assign	SYNTHESIZED_WIRE_170 = B[28] & A[18];

assign	SYNTHESIZED_WIRE_167 = B[28] & A[17];

assign	SYNTHESIZED_WIRE_257 = B[28] & A[16];


OneBitAdder	b2v_inst197(
	.ci(SYNTHESIZED_WIRE_365),
	.a(SYNTHESIZED_WIRE_366),
	.b(SYNTHESIZED_WIRE_367),
	.co(SYNTHESIZED_WIRE_368),
	.s(SYNTHESIZED_WIRE_269));

assign	SYNTHESIZED_WIRE_254 = B[28] & A[15];

assign	SYNTHESIZED_WIRE_251 = B[28] & A[14];

assign	SYNTHESIZED_WIRE_248 = B[28] & A[13];

assign	SYNTHESIZED_WIRE_245 = B[28] & A[12];

assign	SYNTHESIZED_WIRE_242 = B[28] & A[11];

assign	SYNTHESIZED_WIRE_239 = B[28] & A[10];

assign	SYNTHESIZED_WIRE_236 = B[28] & A[9];

assign	SYNTHESIZED_WIRE_233 = B[28] & A[8];

assign	SYNTHESIZED_WIRE_230 = B[28] & A[7];

assign	SYNTHESIZED_WIRE_227 = B[28] & A[6];


OneBitAdder	b2v_inst198(
	.ci(SYNTHESIZED_WIRE_368),
	.a(SYNTHESIZED_WIRE_369),
	.b(SYNTHESIZED_WIRE_370),
	.co(SYNTHESIZED_WIRE_371),
	.s(SYNTHESIZED_WIRE_272));

assign	SYNTHESIZED_WIRE_224 = B[28] & A[5];

assign	SYNTHESIZED_WIRE_221 = B[28] & A[4];

assign	SYNTHESIZED_WIRE_218 = B[28] & A[3];

assign	SYNTHESIZED_WIRE_215 = B[28] & A[2];

assign	SYNTHESIZED_WIRE_212 = B[28] & A[1];

assign	SYNTHESIZED_WIRE_165 = B[28] & A[0];

assign	SYNTHESIZED_WIRE_111 = B[29] & A[30];

assign	SYNTHESIZED_WIRE_114 = ~(A[31] & B[29]);

assign	SYNTHESIZED_WIRE_108 = B[29] & A[29];

assign	SYNTHESIZED_WIRE_105 = B[29] & A[28];


OneBitAdder	b2v_inst199(
	.ci(SYNTHESIZED_WIRE_371),
	.a(SYNTHESIZED_WIRE_372),
	.b(SYNTHESIZED_WIRE_373),
	.co(SYNTHESIZED_WIRE_376),
	.s(SYNTHESIZED_WIRE_275));

assign	SYNTHESIZED_WIRE_102 = B[29] & A[27];

assign	SYNTHESIZED_WIRE_99 = B[29] & A[26];

assign	SYNTHESIZED_WIRE_96 = B[29] & A[25];

assign	SYNTHESIZED_WIRE_93 = B[29] & A[24];

assign	SYNTHESIZED_WIRE_90 = B[29] & A[23];

assign	SYNTHESIZED_WIRE_87 = B[29] & A[22];

assign	SYNTHESIZED_WIRE_69 = B[29] & A[21];

assign	SYNTHESIZED_WIRE_36 = B[29] & A[20];

assign	SYNTHESIZED_WIRE_3 = B[29] & A[19];

assign	SYNTHESIZED_WIRE_2916 = B[29] & A[18];


OneBitAdderHalf	b2v_inst2(
	.A(SYNTHESIZED_WIRE_374),
	.B(SYNTHESIZED_WIRE_375),
	.C(SYNTHESIZED_WIRE_2327),
	.S(Z_ALTERA_SYNTHESIZED[30]));


OneBitAdder	b2v_inst200(
	.ci(SYNTHESIZED_WIRE_376),
	.a(SYNTHESIZED_WIRE_377),
	.b(SYNTHESIZED_WIRE_378),
	.co(SYNTHESIZED_WIRE_379),
	.s(SYNTHESIZED_WIRE_278));

assign	SYNTHESIZED_WIRE_2883 = B[29] & A[17];

assign	SYNTHESIZED_WIRE_162 = B[29] & A[16];

assign	SYNTHESIZED_WIRE_159 = B[29] & A[15];

assign	SYNTHESIZED_WIRE_156 = B[29] & A[14];

assign	SYNTHESIZED_WIRE_153 = B[29] & A[13];

assign	SYNTHESIZED_WIRE_150 = B[29] & A[12];

assign	SYNTHESIZED_WIRE_147 = B[29] & A[11];

assign	SYNTHESIZED_WIRE_144 = B[29] & A[10];

assign	SYNTHESIZED_WIRE_141 = B[29] & A[9];

assign	SYNTHESIZED_WIRE_138 = B[29] & A[8];


OneBitAdder	b2v_inst201(
	.ci(SYNTHESIZED_WIRE_379),
	.a(SYNTHESIZED_WIRE_380),
	.b(SYNTHESIZED_WIRE_381),
	.co(SYNTHESIZED_WIRE_382),
	.s(SYNTHESIZED_WIRE_281));

assign	SYNTHESIZED_WIRE_135 = B[29] & A[7];

assign	SYNTHESIZED_WIRE_132 = B[29] & A[6];

assign	SYNTHESIZED_WIRE_129 = B[29] & A[5];

assign	SYNTHESIZED_WIRE_126 = B[29] & A[4];

assign	SYNTHESIZED_WIRE_123 = B[29] & A[3];

assign	SYNTHESIZED_WIRE_120 = B[29] & A[2];

assign	SYNTHESIZED_WIRE_117 = B[29] & A[1];

assign	SYNTHESIZED_WIRE_2851 = B[29] & A[0];

assign	SYNTHESIZED_WIRE_2263 = B[30] & A[30];

assign	SYNTHESIZED_WIRE_2296 = ~(A[31] & B[30]);


OneBitAdder	b2v_inst202(
	.ci(SYNTHESIZED_WIRE_382),
	.a(SYNTHESIZED_WIRE_383),
	.b(SYNTHESIZED_WIRE_384),
	.co(SYNTHESIZED_WIRE_385),
	.s(SYNTHESIZED_WIRE_284));

assign	SYNTHESIZED_WIRE_2230 = B[30] & A[29];

assign	SYNTHESIZED_WIRE_2197 = B[30] & A[28];

assign	SYNTHESIZED_WIRE_2165 = B[30] & A[27];

assign	SYNTHESIZED_WIRE_2132 = B[30] & A[26];

assign	SYNTHESIZED_WIRE_2099 = B[30] & A[25];

assign	SYNTHESIZED_WIRE_2067 = B[30] & A[24];

assign	SYNTHESIZED_WIRE_2034 = B[30] & A[23];

assign	SYNTHESIZED_WIRE_2001 = B[30] & A[22];

assign	SYNTHESIZED_WIRE_1969 = B[30] & A[21];

assign	SYNTHESIZED_WIRE_1936 = B[30] & A[20];


OneBitAdder	b2v_inst203(
	.ci(SYNTHESIZED_WIRE_385),
	.a(SYNTHESIZED_WIRE_386),
	.b(SYNTHESIZED_WIRE_387),
	.co(SYNTHESIZED_WIRE_388),
	.s(SYNTHESIZED_WIRE_287));

assign	SYNTHESIZED_WIRE_1903 = B[30] & A[19];

assign	SYNTHESIZED_WIRE_1871 = B[30] & A[18];

assign	SYNTHESIZED_WIRE_1838 = B[30] & A[17];

assign	SYNTHESIZED_WIRE_2819 = B[30] & A[16];

assign	SYNTHESIZED_WIRE_2786 = B[30] & A[15];

assign	SYNTHESIZED_WIRE_2753 = B[30] & A[14];

assign	SYNTHESIZED_WIRE_2720 = B[30] & A[13];

assign	SYNTHESIZED_WIRE_2688 = B[30] & A[12];

assign	SYNTHESIZED_WIRE_2655 = B[30] & A[11];

assign	SYNTHESIZED_WIRE_2622 = B[30] & A[10];


OneBitAdder	b2v_inst204(
	.ci(SYNTHESIZED_WIRE_388),
	.a(SYNTHESIZED_WIRE_389),
	.b(SYNTHESIZED_WIRE_390),
	.co(SYNTHESIZED_WIRE_391),
	.s(SYNTHESIZED_WIRE_290));

assign	SYNTHESIZED_WIRE_2590 = B[30] & A[9];

assign	SYNTHESIZED_WIRE_2557 = B[30] & A[8];

assign	SYNTHESIZED_WIRE_2524 = B[30] & A[7];

assign	SYNTHESIZED_WIRE_2492 = B[30] & A[6];

assign	SYNTHESIZED_WIRE_2459 = B[30] & A[5];

assign	SYNTHESIZED_WIRE_2426 = B[30] & A[4];

assign	SYNTHESIZED_WIRE_2394 = B[30] & A[3];

assign	SYNTHESIZED_WIRE_2361 = B[30] & A[2];

assign	SYNTHESIZED_WIRE_2328 = B[30] & A[1];

assign	SYNTHESIZED_WIRE_375 = B[30] & A[0];


OneBitAdder	b2v_inst205(
	.ci(SYNTHESIZED_WIRE_391),
	.a(SYNTHESIZED_WIRE_392),
	.b(SYNTHESIZED_WIRE_393),
	.co(SYNTHESIZED_WIRE_394),
	.s(SYNTHESIZED_WIRE_293));

assign	SYNTHESIZED_WIRE_1315 = ~(A[1] & B[31]);

assign	SYNTHESIZED_WIRE_1348 = ~(A[2] & B[31]);

assign	SYNTHESIZED_WIRE_1380 = ~(A[3] & B[31]);

assign	SYNTHESIZED_WIRE_1413 = ~(A[4] & B[31]);

assign	SYNTHESIZED_WIRE_1446 = ~(A[5] & B[31]);

assign	SYNTHESIZED_WIRE_1478 = ~(A[6] & B[31]);

assign	SYNTHESIZED_WIRE_1511 = ~(A[7] & B[31]);

assign	SYNTHESIZED_WIRE_1544 = ~(A[8] & B[31]);

assign	SYNTHESIZED_WIRE_1576 = ~(A[9] & B[31]);

assign	SYNTHESIZED_WIRE_1609 = ~(A[10] & B[31]);


OneBitAdder	b2v_inst206(
	.ci(SYNTHESIZED_WIRE_394),
	.a(SYNTHESIZED_WIRE_395),
	.b(SYNTHESIZED_WIRE_396),
	.co(SYNTHESIZED_WIRE_397),
	.s(SYNTHESIZED_WIRE_296));

assign	SYNTHESIZED_WIRE_1642 = ~(A[11] & B[31]);

assign	SYNTHESIZED_WIRE_1674 = ~(A[12] & B[31]);

assign	SYNTHESIZED_WIRE_1707 = ~(A[13] & B[31]);

assign	SYNTHESIZED_WIRE_1740 = ~(A[14] & B[31]);

assign	SYNTHESIZED_WIRE_1773 = ~(A[15] & B[31]);

assign	SYNTHESIZED_WIRE_1805 = ~(A[16] & B[31]);

assign	SYNTHESIZED_WIRE_825 = ~(A[17] & B[31]);

assign	SYNTHESIZED_WIRE_857 = ~(A[18] & B[31]);

assign	SYNTHESIZED_WIRE_890 = ~(A[19] & B[31]);

assign	SYNTHESIZED_WIRE_923 = ~(A[20] & B[31]);


OneBitAdder	b2v_inst207(
	.ci(SYNTHESIZED_WIRE_397),
	.a(SYNTHESIZED_WIRE_398),
	.b(SYNTHESIZED_WIRE_399),
	.co(SYNTHESIZED_WIRE_400),
	.s(SYNTHESIZED_WIRE_299));

assign	SYNTHESIZED_WIRE_955 = ~(A[21] & B[31]);

assign	SYNTHESIZED_WIRE_988 = ~(A[22] & B[31]);

assign	SYNTHESIZED_WIRE_1021 = ~(A[23] & B[31]);

assign	SYNTHESIZED_WIRE_1053 = ~(A[24] & B[31]);

assign	SYNTHESIZED_WIRE_1086 = ~(A[25] & B[31]);

assign	SYNTHESIZED_WIRE_1119 = ~(A[26] & B[31]);

assign	SYNTHESIZED_WIRE_1151 = ~(A[27] & B[31]);

assign	SYNTHESIZED_WIRE_1184 = ~(A[28] & B[31]);

assign	SYNTHESIZED_WIRE_1217 = ~(A[29] & B[31]);

assign	SYNTHESIZED_WIRE_1250 = ~(A[30] & B[31]);


OneBitAdder	b2v_inst208(
	.ci(SYNTHESIZED_WIRE_400),
	.a(SYNTHESIZED_WIRE_401),
	.b(SYNTHESIZED_WIRE_402),
	.co(SYNTHESIZED_WIRE_305),
	.s(SYNTHESIZED_WIRE_302));


OneBitAdder	b2v_inst209(
	.ci(SYNTHESIZED_WIRE_403),
	.a(SYNTHESIZED_WIRE_404),
	.b(SYNTHESIZED_WIRE_405),
	.co(SYNTHESIZED_WIRE_406),
	.s(SYNTHESIZED_WIRE_259));


OneBitAdder	b2v_inst210(
	.ci(SYNTHESIZED_WIRE_406),
	.a(SYNTHESIZED_WIRE_407),
	.b(SYNTHESIZED_WIRE_408),
	.co(SYNTHESIZED_WIRE_409),
	.s(SYNTHESIZED_WIRE_308));


OneBitAdder	b2v_inst211(
	.ci(SYNTHESIZED_WIRE_409),
	.a(SYNTHESIZED_WIRE_410),
	.b(SYNTHESIZED_WIRE_411),
	.co(SYNTHESIZED_WIRE_412),
	.s(SYNTHESIZED_WIRE_311));


OneBitAdder	b2v_inst212(
	.ci(SYNTHESIZED_WIRE_412),
	.a(SYNTHESIZED_WIRE_413),
	.b(SYNTHESIZED_WIRE_414),
	.co(SYNTHESIZED_WIRE_415),
	.s(SYNTHESIZED_WIRE_314));


OneBitAdder	b2v_inst213(
	.ci(SYNTHESIZED_WIRE_415),
	.a(SYNTHESIZED_WIRE_416),
	.b(SYNTHESIZED_WIRE_417),
	.co(SYNTHESIZED_WIRE_418),
	.s(SYNTHESIZED_WIRE_317));


OneBitAdder	b2v_inst214(
	.ci(SYNTHESIZED_WIRE_418),
	.a(SYNTHESIZED_WIRE_419),
	.b(SYNTHESIZED_WIRE_420),
	.co(SYNTHESIZED_WIRE_421),
	.s(SYNTHESIZED_WIRE_320));


OneBitAdder	b2v_inst215(
	.ci(SYNTHESIZED_WIRE_421),
	.a(SYNTHESIZED_WIRE_422),
	.b(SYNTHESIZED_WIRE_423),
	.co(SYNTHESIZED_WIRE_424),
	.s(SYNTHESIZED_WIRE_323));


OneBitAdder	b2v_inst216(
	.ci(SYNTHESIZED_WIRE_424),
	.a(SYNTHESIZED_WIRE_425),
	.b(SYNTHESIZED_WIRE_426),
	.co(SYNTHESIZED_WIRE_427),
	.s(SYNTHESIZED_WIRE_326));


OneBitAdder	b2v_inst217(
	.ci(SYNTHESIZED_WIRE_427),
	.a(SYNTHESIZED_WIRE_428),
	.b(SYNTHESIZED_WIRE_429),
	.co(SYNTHESIZED_WIRE_430),
	.s(SYNTHESIZED_WIRE_329));


OneBitAdder	b2v_inst218(
	.ci(SYNTHESIZED_WIRE_430),
	.a(SYNTHESIZED_WIRE_431),
	.b(SYNTHESIZED_WIRE_432),
	.co(SYNTHESIZED_WIRE_433),
	.s(SYNTHESIZED_WIRE_332));


OneBitAdder	b2v_inst219(
	.ci(SYNTHESIZED_WIRE_433),
	.a(SYNTHESIZED_WIRE_434),
	.b(SYNTHESIZED_WIRE_435),
	.co(SYNTHESIZED_WIRE_436),
	.s(SYNTHESIZED_WIRE_335));


OneBitAdder	b2v_inst220(
	.ci(SYNTHESIZED_WIRE_436),
	.a(SYNTHESIZED_WIRE_437),
	.b(SYNTHESIZED_WIRE_438),
	.co(SYNTHESIZED_WIRE_439),
	.s(SYNTHESIZED_WIRE_338));


OneBitAdder	b2v_inst221(
	.ci(SYNTHESIZED_WIRE_439),
	.a(SYNTHESIZED_WIRE_440),
	.b(SYNTHESIZED_WIRE_441),
	.co(SYNTHESIZED_WIRE_442),
	.s(SYNTHESIZED_WIRE_341));


OneBitAdder	b2v_inst222(
	.ci(SYNTHESIZED_WIRE_442),
	.a(SYNTHESIZED_WIRE_443),
	.b(SYNTHESIZED_WIRE_444),
	.co(SYNTHESIZED_WIRE_445),
	.s(SYNTHESIZED_WIRE_344));


OneBitAdder	b2v_inst223(
	.ci(SYNTHESIZED_WIRE_445),
	.a(SYNTHESIZED_WIRE_446),
	.b(SYNTHESIZED_WIRE_447),
	.co(SYNTHESIZED_WIRE_448),
	.s(SYNTHESIZED_WIRE_347));


OneBitAdder	b2v_inst224(
	.ci(SYNTHESIZED_WIRE_448),
	.a(SYNTHESIZED_WIRE_449),
	.b(SYNTHESIZED_WIRE_450),
	.co(SYNTHESIZED_WIRE_356),
	.s(SYNTHESIZED_WIRE_350));


OneBitAdderHalf	b2v_inst225(
	.A(SYNTHESIZED_WIRE_451),
	.B(SYNTHESIZED_WIRE_452),
	.C(SYNTHESIZED_WIRE_498),
	.S(Z_ALTERA_SYNTHESIZED[25]));


OneBitAdder	b2v_inst226(
	.ci(SYNTHESIZED_WIRE_453),
	.a(SYNTHESIZED_WIRE_454),
	.b(SYNTHESIZED_WIRE_455),
	.co(SYNTHESIZED_WIRE_456),
	.s(SYNTHESIZED_WIRE_450));


OneBitAdder	b2v_inst227(
	.ci(SYNTHESIZED_WIRE_456),
	.a(SYNTHESIZED_WIRE_457),
	.b(SYNTHESIZED_WIRE_458),
	.co(SYNTHESIZED_WIRE_459),
	.s(SYNTHESIZED_WIRE_358));


OneBitAdder	b2v_inst228(
	.ci(SYNTHESIZED_WIRE_459),
	.a(SYNTHESIZED_WIRE_460),
	.b(SYNTHESIZED_WIRE_461),
	.co(SYNTHESIZED_WIRE_462),
	.s(SYNTHESIZED_WIRE_361));


OneBitAdder	b2v_inst229(
	.ci(SYNTHESIZED_WIRE_462),
	.a(SYNTHESIZED_WIRE_463),
	.b(SYNTHESIZED_WIRE_464),
	.co(SYNTHESIZED_WIRE_465),
	.s(SYNTHESIZED_WIRE_364));


OneBitAdder	b2v_inst230(
	.ci(SYNTHESIZED_WIRE_465),
	.a(SYNTHESIZED_WIRE_466),
	.b(SYNTHESIZED_WIRE_467),
	.co(SYNTHESIZED_WIRE_468),
	.s(SYNTHESIZED_WIRE_367));


OneBitAdder	b2v_inst231(
	.ci(SYNTHESIZED_WIRE_468),
	.a(SYNTHESIZED_WIRE_469),
	.b(SYNTHESIZED_WIRE_470),
	.co(SYNTHESIZED_WIRE_471),
	.s(SYNTHESIZED_WIRE_370));


OneBitAdder	b2v_inst232(
	.ci(SYNTHESIZED_WIRE_471),
	.a(SYNTHESIZED_WIRE_472),
	.b(SYNTHESIZED_WIRE_473),
	.co(SYNTHESIZED_WIRE_474),
	.s(SYNTHESIZED_WIRE_373));


OneBitAdder	b2v_inst233(
	.ci(SYNTHESIZED_WIRE_474),
	.a(SYNTHESIZED_WIRE_475),
	.b(SYNTHESIZED_WIRE_476),
	.co(SYNTHESIZED_WIRE_477),
	.s(SYNTHESIZED_WIRE_378));


OneBitAdder	b2v_inst234(
	.ci(SYNTHESIZED_WIRE_477),
	.a(SYNTHESIZED_WIRE_478),
	.b(SYNTHESIZED_WIRE_479),
	.co(SYNTHESIZED_WIRE_480),
	.s(SYNTHESIZED_WIRE_381));


OneBitAdder	b2v_inst235(
	.ci(SYNTHESIZED_WIRE_480),
	.a(SYNTHESIZED_WIRE_481),
	.b(SYNTHESIZED_WIRE_482),
	.co(SYNTHESIZED_WIRE_483),
	.s(SYNTHESIZED_WIRE_384));


OneBitAdder	b2v_inst236(
	.ci(SYNTHESIZED_WIRE_483),
	.a(SYNTHESIZED_WIRE_484),
	.b(SYNTHESIZED_WIRE_485),
	.co(SYNTHESIZED_WIRE_486),
	.s(SYNTHESIZED_WIRE_387));


OneBitAdder	b2v_inst237(
	.ci(SYNTHESIZED_WIRE_486),
	.a(SYNTHESIZED_WIRE_487),
	.b(SYNTHESIZED_WIRE_488),
	.co(SYNTHESIZED_WIRE_489),
	.s(SYNTHESIZED_WIRE_390));


OneBitAdder	b2v_inst238(
	.ci(SYNTHESIZED_WIRE_489),
	.a(SYNTHESIZED_WIRE_490),
	.b(SYNTHESIZED_WIRE_491),
	.co(SYNTHESIZED_WIRE_492),
	.s(SYNTHESIZED_WIRE_393));


OneBitAdder	b2v_inst239(
	.ci(SYNTHESIZED_WIRE_492),
	.a(SYNTHESIZED_WIRE_493),
	.b(SYNTHESIZED_WIRE_494),
	.co(SYNTHESIZED_WIRE_495),
	.s(SYNTHESIZED_WIRE_396));


OneBitAdder	b2v_inst240(
	.ci(SYNTHESIZED_WIRE_495),
	.a(SYNTHESIZED_WIRE_496),
	.b(SYNTHESIZED_WIRE_497),
	.co(SYNTHESIZED_WIRE_402),
	.s(SYNTHESIZED_WIRE_399));


OneBitAdder	b2v_inst241(
	.ci(SYNTHESIZED_WIRE_498),
	.a(SYNTHESIZED_WIRE_499),
	.b(SYNTHESIZED_WIRE_500),
	.co(SYNTHESIZED_WIRE_501),
	.s(SYNTHESIZED_WIRE_354));


OneBitAdder	b2v_inst242(
	.ci(SYNTHESIZED_WIRE_501),
	.a(SYNTHESIZED_WIRE_502),
	.b(SYNTHESIZED_WIRE_503),
	.co(SYNTHESIZED_WIRE_504),
	.s(SYNTHESIZED_WIRE_405));


OneBitAdder	b2v_inst243(
	.ci(SYNTHESIZED_WIRE_504),
	.a(SYNTHESIZED_WIRE_505),
	.b(SYNTHESIZED_WIRE_506),
	.co(SYNTHESIZED_WIRE_507),
	.s(SYNTHESIZED_WIRE_408));


OneBitAdder	b2v_inst244(
	.ci(SYNTHESIZED_WIRE_507),
	.a(SYNTHESIZED_WIRE_508),
	.b(SYNTHESIZED_WIRE_509),
	.co(SYNTHESIZED_WIRE_510),
	.s(SYNTHESIZED_WIRE_411));


OneBitAdder	b2v_inst245(
	.ci(SYNTHESIZED_WIRE_510),
	.a(SYNTHESIZED_WIRE_511),
	.b(SYNTHESIZED_WIRE_512),
	.co(SYNTHESIZED_WIRE_513),
	.s(SYNTHESIZED_WIRE_414));


OneBitAdder	b2v_inst246(
	.ci(SYNTHESIZED_WIRE_513),
	.a(SYNTHESIZED_WIRE_514),
	.b(SYNTHESIZED_WIRE_515),
	.co(SYNTHESIZED_WIRE_516),
	.s(SYNTHESIZED_WIRE_417));


OneBitAdder	b2v_inst247(
	.ci(SYNTHESIZED_WIRE_516),
	.a(SYNTHESIZED_WIRE_517),
	.b(SYNTHESIZED_WIRE_518),
	.co(SYNTHESIZED_WIRE_519),
	.s(SYNTHESIZED_WIRE_420));


OneBitAdder	b2v_inst248(
	.ci(SYNTHESIZED_WIRE_519),
	.a(SYNTHESIZED_WIRE_520),
	.b(SYNTHESIZED_WIRE_521),
	.co(SYNTHESIZED_WIRE_522),
	.s(SYNTHESIZED_WIRE_423));


OneBitAdder	b2v_inst249(
	.ci(SYNTHESIZED_WIRE_522),
	.a(SYNTHESIZED_WIRE_523),
	.b(SYNTHESIZED_WIRE_524),
	.co(SYNTHESIZED_WIRE_525),
	.s(SYNTHESIZED_WIRE_426));


OneBitAdder	b2v_inst250(
	.ci(SYNTHESIZED_WIRE_525),
	.a(SYNTHESIZED_WIRE_526),
	.b(SYNTHESIZED_WIRE_527),
	.co(SYNTHESIZED_WIRE_528),
	.s(SYNTHESIZED_WIRE_429));


OneBitAdder	b2v_inst251(
	.ci(SYNTHESIZED_WIRE_528),
	.a(SYNTHESIZED_WIRE_529),
	.b(SYNTHESIZED_WIRE_530),
	.co(SYNTHESIZED_WIRE_531),
	.s(SYNTHESIZED_WIRE_432));


OneBitAdder	b2v_inst252(
	.ci(SYNTHESIZED_WIRE_531),
	.a(SYNTHESIZED_WIRE_532),
	.b(SYNTHESIZED_WIRE_533),
	.co(SYNTHESIZED_WIRE_534),
	.s(SYNTHESIZED_WIRE_435));


OneBitAdder	b2v_inst253(
	.ci(SYNTHESIZED_WIRE_534),
	.a(SYNTHESIZED_WIRE_535),
	.b(SYNTHESIZED_WIRE_536),
	.co(SYNTHESIZED_WIRE_537),
	.s(SYNTHESIZED_WIRE_438));


OneBitAdder	b2v_inst254(
	.ci(SYNTHESIZED_WIRE_537),
	.a(SYNTHESIZED_WIRE_538),
	.b(SYNTHESIZED_WIRE_539),
	.co(SYNTHESIZED_WIRE_540),
	.s(SYNTHESIZED_WIRE_441));


OneBitAdder	b2v_inst255(
	.ci(SYNTHESIZED_WIRE_540),
	.a(SYNTHESIZED_WIRE_541),
	.b(SYNTHESIZED_WIRE_542),
	.co(SYNTHESIZED_WIRE_543),
	.s(SYNTHESIZED_WIRE_444));


OneBitAdder	b2v_inst256(
	.ci(SYNTHESIZED_WIRE_543),
	.a(SYNTHESIZED_WIRE_544),
	.b(SYNTHESIZED_WIRE_545),
	.co(SYNTHESIZED_WIRE_453),
	.s(SYNTHESIZED_WIRE_447));


OneBitAdderHalf	b2v_inst257(
	.A(SYNTHESIZED_WIRE_546),
	.B(SYNTHESIZED_WIRE_547),
	.C(SYNTHESIZED_WIRE_593),
	.S(Z_ALTERA_SYNTHESIZED[24]));


OneBitAdder	b2v_inst258(
	.ci(SYNTHESIZED_WIRE_548),
	.a(SYNTHESIZED_WIRE_549),
	.b(SYNTHESIZED_WIRE_550),
	.co(SYNTHESIZED_WIRE_551),
	.s(SYNTHESIZED_WIRE_545));


OneBitAdder	b2v_inst259(
	.ci(SYNTHESIZED_WIRE_551),
	.a(SYNTHESIZED_WIRE_552),
	.b(SYNTHESIZED_WIRE_553),
	.co(SYNTHESIZED_WIRE_554),
	.s(SYNTHESIZED_WIRE_455));


OneBitAdder	b2v_inst260(
	.ci(SYNTHESIZED_WIRE_554),
	.a(SYNTHESIZED_WIRE_555),
	.b(SYNTHESIZED_WIRE_556),
	.co(SYNTHESIZED_WIRE_557),
	.s(SYNTHESIZED_WIRE_458));


OneBitAdder	b2v_inst261(
	.ci(SYNTHESIZED_WIRE_557),
	.a(SYNTHESIZED_WIRE_558),
	.b(SYNTHESIZED_WIRE_559),
	.co(SYNTHESIZED_WIRE_560),
	.s(SYNTHESIZED_WIRE_461));


OneBitAdder	b2v_inst262(
	.ci(SYNTHESIZED_WIRE_560),
	.a(SYNTHESIZED_WIRE_561),
	.b(SYNTHESIZED_WIRE_562),
	.co(SYNTHESIZED_WIRE_563),
	.s(SYNTHESIZED_WIRE_464));


OneBitAdder	b2v_inst263(
	.ci(SYNTHESIZED_WIRE_563),
	.a(SYNTHESIZED_WIRE_564),
	.b(SYNTHESIZED_WIRE_565),
	.co(SYNTHESIZED_WIRE_566),
	.s(SYNTHESIZED_WIRE_467));


OneBitAdder	b2v_inst264(
	.ci(SYNTHESIZED_WIRE_566),
	.a(SYNTHESIZED_WIRE_567),
	.b(SYNTHESIZED_WIRE_568),
	.co(SYNTHESIZED_WIRE_569),
	.s(SYNTHESIZED_WIRE_470));


OneBitAdder	b2v_inst265(
	.ci(SYNTHESIZED_WIRE_569),
	.a(SYNTHESIZED_WIRE_570),
	.b(SYNTHESIZED_WIRE_571),
	.co(SYNTHESIZED_WIRE_572),
	.s(SYNTHESIZED_WIRE_473));


OneBitAdder	b2v_inst266(
	.ci(SYNTHESIZED_WIRE_572),
	.a(SYNTHESIZED_WIRE_573),
	.b(SYNTHESIZED_WIRE_574),
	.co(SYNTHESIZED_WIRE_575),
	.s(SYNTHESIZED_WIRE_476));


OneBitAdder	b2v_inst267(
	.ci(SYNTHESIZED_WIRE_575),
	.a(SYNTHESIZED_WIRE_576),
	.b(SYNTHESIZED_WIRE_577),
	.co(SYNTHESIZED_WIRE_578),
	.s(SYNTHESIZED_WIRE_479));


OneBitAdder	b2v_inst268(
	.ci(SYNTHESIZED_WIRE_578),
	.a(SYNTHESIZED_WIRE_579),
	.b(SYNTHESIZED_WIRE_580),
	.co(SYNTHESIZED_WIRE_581),
	.s(SYNTHESIZED_WIRE_482));


OneBitAdder	b2v_inst269(
	.ci(SYNTHESIZED_WIRE_581),
	.a(SYNTHESIZED_WIRE_582),
	.b(SYNTHESIZED_WIRE_583),
	.co(SYNTHESIZED_WIRE_584),
	.s(SYNTHESIZED_WIRE_485));


OneBitAdder	b2v_inst270(
	.ci(SYNTHESIZED_WIRE_584),
	.a(SYNTHESIZED_WIRE_585),
	.b(SYNTHESIZED_WIRE_586),
	.co(SYNTHESIZED_WIRE_587),
	.s(SYNTHESIZED_WIRE_488));


OneBitAdder	b2v_inst271(
	.ci(SYNTHESIZED_WIRE_587),
	.a(SYNTHESIZED_WIRE_588),
	.b(SYNTHESIZED_WIRE_589),
	.co(SYNTHESIZED_WIRE_590),
	.s(SYNTHESIZED_WIRE_491));


OneBitAdder	b2v_inst272(
	.ci(SYNTHESIZED_WIRE_590),
	.a(SYNTHESIZED_WIRE_591),
	.b(SYNTHESIZED_WIRE_592),
	.co(SYNTHESIZED_WIRE_497),
	.s(SYNTHESIZED_WIRE_494));


OneBitAdder	b2v_inst273(
	.ci(SYNTHESIZED_WIRE_593),
	.a(SYNTHESIZED_WIRE_594),
	.b(SYNTHESIZED_WIRE_595),
	.co(SYNTHESIZED_WIRE_596),
	.s(SYNTHESIZED_WIRE_451));


OneBitAdder	b2v_inst274(
	.ci(SYNTHESIZED_WIRE_596),
	.a(SYNTHESIZED_WIRE_597),
	.b(SYNTHESIZED_WIRE_598),
	.co(SYNTHESIZED_WIRE_599),
	.s(SYNTHESIZED_WIRE_500));


OneBitAdder	b2v_inst275(
	.ci(SYNTHESIZED_WIRE_599),
	.a(SYNTHESIZED_WIRE_600),
	.b(SYNTHESIZED_WIRE_601),
	.co(SYNTHESIZED_WIRE_602),
	.s(SYNTHESIZED_WIRE_503));


OneBitAdder	b2v_inst276(
	.ci(SYNTHESIZED_WIRE_602),
	.a(SYNTHESIZED_WIRE_603),
	.b(SYNTHESIZED_WIRE_604),
	.co(SYNTHESIZED_WIRE_605),
	.s(SYNTHESIZED_WIRE_506));


OneBitAdder	b2v_inst277(
	.ci(SYNTHESIZED_WIRE_605),
	.a(SYNTHESIZED_WIRE_606),
	.b(SYNTHESIZED_WIRE_607),
	.co(SYNTHESIZED_WIRE_608),
	.s(SYNTHESIZED_WIRE_509));


OneBitAdder	b2v_inst278(
	.ci(SYNTHESIZED_WIRE_608),
	.a(SYNTHESIZED_WIRE_609),
	.b(SYNTHESIZED_WIRE_610),
	.co(SYNTHESIZED_WIRE_611),
	.s(SYNTHESIZED_WIRE_512));


OneBitAdder	b2v_inst279(
	.ci(SYNTHESIZED_WIRE_611),
	.a(SYNTHESIZED_WIRE_612),
	.b(SYNTHESIZED_WIRE_613),
	.co(SYNTHESIZED_WIRE_614),
	.s(SYNTHESIZED_WIRE_515));


OneBitAdder	b2v_inst280(
	.ci(SYNTHESIZED_WIRE_614),
	.a(SYNTHESIZED_WIRE_615),
	.b(SYNTHESIZED_WIRE_616),
	.co(SYNTHESIZED_WIRE_617),
	.s(SYNTHESIZED_WIRE_518));


OneBitAdder	b2v_inst281(
	.ci(SYNTHESIZED_WIRE_617),
	.a(SYNTHESIZED_WIRE_618),
	.b(SYNTHESIZED_WIRE_619),
	.co(SYNTHESIZED_WIRE_620),
	.s(SYNTHESIZED_WIRE_521));


OneBitAdder	b2v_inst282(
	.ci(SYNTHESIZED_WIRE_620),
	.a(SYNTHESIZED_WIRE_621),
	.b(SYNTHESIZED_WIRE_622),
	.co(SYNTHESIZED_WIRE_623),
	.s(SYNTHESIZED_WIRE_524));


OneBitAdder	b2v_inst283(
	.ci(SYNTHESIZED_WIRE_623),
	.a(SYNTHESIZED_WIRE_624),
	.b(SYNTHESIZED_WIRE_625),
	.co(SYNTHESIZED_WIRE_626),
	.s(SYNTHESIZED_WIRE_527));


OneBitAdder	b2v_inst284(
	.ci(SYNTHESIZED_WIRE_626),
	.a(SYNTHESIZED_WIRE_627),
	.b(SYNTHESIZED_WIRE_628),
	.co(SYNTHESIZED_WIRE_629),
	.s(SYNTHESIZED_WIRE_530));


OneBitAdder	b2v_inst285(
	.ci(SYNTHESIZED_WIRE_629),
	.a(SYNTHESIZED_WIRE_630),
	.b(SYNTHESIZED_WIRE_631),
	.co(SYNTHESIZED_WIRE_632),
	.s(SYNTHESIZED_WIRE_533));


OneBitAdder	b2v_inst286(
	.ci(SYNTHESIZED_WIRE_632),
	.a(SYNTHESIZED_WIRE_633),
	.b(SYNTHESIZED_WIRE_634),
	.co(SYNTHESIZED_WIRE_635),
	.s(SYNTHESIZED_WIRE_536));


OneBitAdder	b2v_inst287(
	.ci(SYNTHESIZED_WIRE_635),
	.a(SYNTHESIZED_WIRE_636),
	.b(SYNTHESIZED_WIRE_637),
	.co(SYNTHESIZED_WIRE_638),
	.s(SYNTHESIZED_WIRE_539));


OneBitAdder	b2v_inst288(
	.ci(SYNTHESIZED_WIRE_638),
	.a(SYNTHESIZED_WIRE_639),
	.b(SYNTHESIZED_WIRE_640),
	.co(SYNTHESIZED_WIRE_548),
	.s(SYNTHESIZED_WIRE_542));


OneBitAdderHalf	b2v_inst289(
	.A(SYNTHESIZED_WIRE_641),
	.B(SYNTHESIZED_WIRE_642),
	.C(SYNTHESIZED_WIRE_690),
	.S(Z_ALTERA_SYNTHESIZED[23]));


OneBitAdder	b2v_inst290(
	.ci(SYNTHESIZED_WIRE_643),
	.a(SYNTHESIZED_WIRE_644),
	.b(SYNTHESIZED_WIRE_645),
	.co(SYNTHESIZED_WIRE_646),
	.s(SYNTHESIZED_WIRE_640));


OneBitAdder	b2v_inst291(
	.ci(SYNTHESIZED_WIRE_646),
	.a(SYNTHESIZED_WIRE_647),
	.b(SYNTHESIZED_WIRE_648),
	.co(SYNTHESIZED_WIRE_649),
	.s(SYNTHESIZED_WIRE_550));


OneBitAdder	b2v_inst292(
	.ci(SYNTHESIZED_WIRE_649),
	.a(SYNTHESIZED_WIRE_650),
	.b(SYNTHESIZED_WIRE_651),
	.co(SYNTHESIZED_WIRE_652),
	.s(SYNTHESIZED_WIRE_553));


OneBitAdder	b2v_inst293(
	.ci(SYNTHESIZED_WIRE_652),
	.a(SYNTHESIZED_WIRE_653),
	.b(SYNTHESIZED_WIRE_654),
	.co(SYNTHESIZED_WIRE_655),
	.s(SYNTHESIZED_WIRE_556));


OneBitAdder	b2v_inst294(
	.ci(SYNTHESIZED_WIRE_655),
	.a(SYNTHESIZED_WIRE_656),
	.b(SYNTHESIZED_WIRE_657),
	.co(SYNTHESIZED_WIRE_658),
	.s(SYNTHESIZED_WIRE_559));


OneBitAdder	b2v_inst295(
	.ci(SYNTHESIZED_WIRE_658),
	.a(SYNTHESIZED_WIRE_659),
	.b(SYNTHESIZED_WIRE_660),
	.co(SYNTHESIZED_WIRE_661),
	.s(SYNTHESIZED_WIRE_562));


OneBitAdder	b2v_inst296(
	.ci(SYNTHESIZED_WIRE_661),
	.a(SYNTHESIZED_WIRE_662),
	.b(SYNTHESIZED_WIRE_663),
	.co(SYNTHESIZED_WIRE_664),
	.s(SYNTHESIZED_WIRE_565));


OneBitAdder	b2v_inst297(
	.ci(SYNTHESIZED_WIRE_664),
	.a(SYNTHESIZED_WIRE_665),
	.b(SYNTHESIZED_WIRE_666),
	.co(SYNTHESIZED_WIRE_667),
	.s(SYNTHESIZED_WIRE_568));


OneBitAdder	b2v_inst298(
	.ci(SYNTHESIZED_WIRE_667),
	.a(SYNTHESIZED_WIRE_668),
	.b(SYNTHESIZED_WIRE_669),
	.co(SYNTHESIZED_WIRE_670),
	.s(SYNTHESIZED_WIRE_571));


OneBitAdder	b2v_inst299(
	.ci(SYNTHESIZED_WIRE_670),
	.a(SYNTHESIZED_WIRE_671),
	.b(SYNTHESIZED_WIRE_672),
	.co(SYNTHESIZED_WIRE_675),
	.s(SYNTHESIZED_WIRE_574));


OneBitAdderHalf	b2v_inst3(
	.A(SYNTHESIZED_WIRE_673),
	.B(SYNTHESIZED_WIRE_674),
	
	.S(Z_ALTERA_SYNTHESIZED[63]));


OneBitAdder	b2v_inst300(
	.ci(SYNTHESIZED_WIRE_675),
	.a(SYNTHESIZED_WIRE_676),
	.b(SYNTHESIZED_WIRE_677),
	.co(SYNTHESIZED_WIRE_678),
	.s(SYNTHESIZED_WIRE_577));


OneBitAdder	b2v_inst301(
	.ci(SYNTHESIZED_WIRE_678),
	.a(SYNTHESIZED_WIRE_679),
	.b(SYNTHESIZED_WIRE_680),
	.co(SYNTHESIZED_WIRE_681),
	.s(SYNTHESIZED_WIRE_580));


OneBitAdder	b2v_inst302(
	.ci(SYNTHESIZED_WIRE_681),
	.a(SYNTHESIZED_WIRE_682),
	.b(SYNTHESIZED_WIRE_683),
	.co(SYNTHESIZED_WIRE_684),
	.s(SYNTHESIZED_WIRE_583));


OneBitAdder	b2v_inst303(
	.ci(SYNTHESIZED_WIRE_684),
	.a(SYNTHESIZED_WIRE_685),
	.b(SYNTHESIZED_WIRE_686),
	.co(SYNTHESIZED_WIRE_687),
	.s(SYNTHESIZED_WIRE_586));


OneBitAdder	b2v_inst304(
	.ci(SYNTHESIZED_WIRE_687),
	.a(SYNTHESIZED_WIRE_688),
	.b(SYNTHESIZED_WIRE_689),
	.co(SYNTHESIZED_WIRE_592),
	.s(SYNTHESIZED_WIRE_589));


OneBitAdder	b2v_inst305(
	.ci(SYNTHESIZED_WIRE_690),
	.a(SYNTHESIZED_WIRE_691),
	.b(SYNTHESIZED_WIRE_692),
	.co(SYNTHESIZED_WIRE_693),
	.s(SYNTHESIZED_WIRE_546));


OneBitAdder	b2v_inst306(
	.ci(SYNTHESIZED_WIRE_693),
	.a(SYNTHESIZED_WIRE_694),
	.b(SYNTHESIZED_WIRE_695),
	.co(SYNTHESIZED_WIRE_696),
	.s(SYNTHESIZED_WIRE_595));


OneBitAdder	b2v_inst307(
	.ci(SYNTHESIZED_WIRE_696),
	.a(SYNTHESIZED_WIRE_697),
	.b(SYNTHESIZED_WIRE_698),
	.co(SYNTHESIZED_WIRE_699),
	.s(SYNTHESIZED_WIRE_598));


OneBitAdder	b2v_inst308(
	.ci(SYNTHESIZED_WIRE_699),
	.a(SYNTHESIZED_WIRE_700),
	.b(SYNTHESIZED_WIRE_701),
	.co(SYNTHESIZED_WIRE_702),
	.s(SYNTHESIZED_WIRE_601));


OneBitAdder	b2v_inst309(
	.ci(SYNTHESIZED_WIRE_702),
	.a(SYNTHESIZED_WIRE_703),
	.b(SYNTHESIZED_WIRE_704),
	.co(SYNTHESIZED_WIRE_705),
	.s(SYNTHESIZED_WIRE_604));


OneBitAdder	b2v_inst310(
	.ci(SYNTHESIZED_WIRE_705),
	.a(SYNTHESIZED_WIRE_706),
	.b(SYNTHESIZED_WIRE_707),
	.co(SYNTHESIZED_WIRE_708),
	.s(SYNTHESIZED_WIRE_607));


OneBitAdder	b2v_inst311(
	.ci(SYNTHESIZED_WIRE_708),
	.a(SYNTHESIZED_WIRE_709),
	.b(SYNTHESIZED_WIRE_710),
	.co(SYNTHESIZED_WIRE_711),
	.s(SYNTHESIZED_WIRE_610));


OneBitAdder	b2v_inst312(
	.ci(SYNTHESIZED_WIRE_711),
	.a(SYNTHESIZED_WIRE_712),
	.b(SYNTHESIZED_WIRE_713),
	.co(SYNTHESIZED_WIRE_714),
	.s(SYNTHESIZED_WIRE_613));


OneBitAdder	b2v_inst313(
	.ci(SYNTHESIZED_WIRE_714),
	.a(SYNTHESIZED_WIRE_715),
	.b(SYNTHESIZED_WIRE_716),
	.co(SYNTHESIZED_WIRE_717),
	.s(SYNTHESIZED_WIRE_616));


OneBitAdder	b2v_inst314(
	.ci(SYNTHESIZED_WIRE_717),
	.a(SYNTHESIZED_WIRE_718),
	.b(SYNTHESIZED_WIRE_719),
	.co(SYNTHESIZED_WIRE_720),
	.s(SYNTHESIZED_WIRE_619));


OneBitAdder	b2v_inst315(
	.ci(SYNTHESIZED_WIRE_720),
	.a(SYNTHESIZED_WIRE_721),
	.b(SYNTHESIZED_WIRE_722),
	.co(SYNTHESIZED_WIRE_723),
	.s(SYNTHESIZED_WIRE_622));


OneBitAdder	b2v_inst316(
	.ci(SYNTHESIZED_WIRE_723),
	.a(SYNTHESIZED_WIRE_724),
	.b(SYNTHESIZED_WIRE_725),
	.co(SYNTHESIZED_WIRE_726),
	.s(SYNTHESIZED_WIRE_625));


OneBitAdder	b2v_inst317(
	.ci(SYNTHESIZED_WIRE_726),
	.a(SYNTHESIZED_WIRE_727),
	.b(SYNTHESIZED_WIRE_728),
	.co(SYNTHESIZED_WIRE_729),
	.s(SYNTHESIZED_WIRE_628));


OneBitAdder	b2v_inst318(
	.ci(SYNTHESIZED_WIRE_729),
	.a(SYNTHESIZED_WIRE_730),
	.b(SYNTHESIZED_WIRE_731),
	.co(SYNTHESIZED_WIRE_732),
	.s(SYNTHESIZED_WIRE_631));


OneBitAdder	b2v_inst319(
	.ci(SYNTHESIZED_WIRE_732),
	.a(SYNTHESIZED_WIRE_733),
	.b(SYNTHESIZED_WIRE_734),
	.co(SYNTHESIZED_WIRE_735),
	.s(SYNTHESIZED_WIRE_634));


OneBitAdder	b2v_inst320(
	.ci(SYNTHESIZED_WIRE_735),
	.a(SYNTHESIZED_WIRE_736),
	.b(SYNTHESIZED_WIRE_737),
	.co(SYNTHESIZED_WIRE_643),
	.s(SYNTHESIZED_WIRE_637));


OneBitAdderHalf	b2v_inst321(
	.A(SYNTHESIZED_WIRE_738),
	.B(SYNTHESIZED_WIRE_739),
	.C(SYNTHESIZED_WIRE_785),
	.S(Z_ALTERA_SYNTHESIZED[22]));


OneBitAdder	b2v_inst322(
	.ci(SYNTHESIZED_WIRE_740),
	.a(SYNTHESIZED_WIRE_741),
	.b(SYNTHESIZED_WIRE_742),
	.co(SYNTHESIZED_WIRE_743),
	.s(SYNTHESIZED_WIRE_737));


OneBitAdder	b2v_inst323(
	.ci(SYNTHESIZED_WIRE_743),
	.a(SYNTHESIZED_WIRE_744),
	.b(SYNTHESIZED_WIRE_745),
	.co(SYNTHESIZED_WIRE_746),
	.s(SYNTHESIZED_WIRE_645));


OneBitAdder	b2v_inst324(
	.ci(SYNTHESIZED_WIRE_746),
	.a(SYNTHESIZED_WIRE_747),
	.b(SYNTHESIZED_WIRE_748),
	.co(SYNTHESIZED_WIRE_749),
	.s(SYNTHESIZED_WIRE_648));


OneBitAdder	b2v_inst325(
	.ci(SYNTHESIZED_WIRE_749),
	.a(SYNTHESIZED_WIRE_750),
	.b(SYNTHESIZED_WIRE_751),
	.co(SYNTHESIZED_WIRE_752),
	.s(SYNTHESIZED_WIRE_651));


OneBitAdder	b2v_inst326(
	.ci(SYNTHESIZED_WIRE_752),
	.a(SYNTHESIZED_WIRE_753),
	.b(SYNTHESIZED_WIRE_754),
	.co(SYNTHESIZED_WIRE_755),
	.s(SYNTHESIZED_WIRE_654));


OneBitAdder	b2v_inst327(
	.ci(SYNTHESIZED_WIRE_755),
	.a(SYNTHESIZED_WIRE_756),
	.b(SYNTHESIZED_WIRE_757),
	.co(SYNTHESIZED_WIRE_758),
	.s(SYNTHESIZED_WIRE_657));


OneBitAdder	b2v_inst328(
	.ci(SYNTHESIZED_WIRE_758),
	.a(SYNTHESIZED_WIRE_759),
	.b(SYNTHESIZED_WIRE_760),
	.co(SYNTHESIZED_WIRE_761),
	.s(SYNTHESIZED_WIRE_660));


OneBitAdder	b2v_inst329(
	.ci(SYNTHESIZED_WIRE_761),
	.a(SYNTHESIZED_WIRE_762),
	.b(SYNTHESIZED_WIRE_763),
	.co(SYNTHESIZED_WIRE_764),
	.s(SYNTHESIZED_WIRE_663));


OneBitAdder	b2v_inst330(
	.ci(SYNTHESIZED_WIRE_764),
	.a(SYNTHESIZED_WIRE_765),
	.b(SYNTHESIZED_WIRE_766),
	.co(SYNTHESIZED_WIRE_767),
	.s(SYNTHESIZED_WIRE_666));


OneBitAdder	b2v_inst331(
	.ci(SYNTHESIZED_WIRE_767),
	.a(SYNTHESIZED_WIRE_768),
	.b(SYNTHESIZED_WIRE_769),
	.co(SYNTHESIZED_WIRE_770),
	.s(SYNTHESIZED_WIRE_669));


OneBitAdder	b2v_inst332(
	.ci(SYNTHESIZED_WIRE_770),
	.a(SYNTHESIZED_WIRE_771),
	.b(SYNTHESIZED_WIRE_772),
	.co(SYNTHESIZED_WIRE_773),
	.s(SYNTHESIZED_WIRE_672));


OneBitAdder	b2v_inst333(
	.ci(SYNTHESIZED_WIRE_773),
	.a(SYNTHESIZED_WIRE_774),
	.b(SYNTHESIZED_WIRE_775),
	.co(SYNTHESIZED_WIRE_776),
	.s(SYNTHESIZED_WIRE_677));


OneBitAdder	b2v_inst334(
	.ci(SYNTHESIZED_WIRE_776),
	.a(SYNTHESIZED_WIRE_777),
	.b(SYNTHESIZED_WIRE_778),
	.co(SYNTHESIZED_WIRE_779),
	.s(SYNTHESIZED_WIRE_680));


OneBitAdder	b2v_inst335(
	.ci(SYNTHESIZED_WIRE_779),
	.a(SYNTHESIZED_WIRE_780),
	.b(SYNTHESIZED_WIRE_781),
	.co(SYNTHESIZED_WIRE_782),
	.s(SYNTHESIZED_WIRE_683));


OneBitAdder	b2v_inst336(
	.ci(SYNTHESIZED_WIRE_782),
	.a(SYNTHESIZED_WIRE_783),
	.b(SYNTHESIZED_WIRE_784),
	.co(SYNTHESIZED_WIRE_689),
	.s(SYNTHESIZED_WIRE_686));


OneBitAdder	b2v_inst337(
	.ci(SYNTHESIZED_WIRE_785),
	.a(SYNTHESIZED_WIRE_786),
	.b(SYNTHESIZED_WIRE_787),
	.co(SYNTHESIZED_WIRE_788),
	.s(SYNTHESIZED_WIRE_641));


OneBitAdder	b2v_inst338(
	.ci(SYNTHESIZED_WIRE_788),
	.a(SYNTHESIZED_WIRE_789),
	.b(SYNTHESIZED_WIRE_790),
	.co(SYNTHESIZED_WIRE_791),
	.s(SYNTHESIZED_WIRE_692));


OneBitAdder	b2v_inst339(
	.ci(SYNTHESIZED_WIRE_791),
	.a(SYNTHESIZED_WIRE_792),
	.b(SYNTHESIZED_WIRE_793),
	.co(SYNTHESIZED_WIRE_794),
	.s(SYNTHESIZED_WIRE_695));


OneBitAdder	b2v_inst340(
	.ci(SYNTHESIZED_WIRE_794),
	.a(SYNTHESIZED_WIRE_795),
	.b(SYNTHESIZED_WIRE_796),
	.co(SYNTHESIZED_WIRE_797),
	.s(SYNTHESIZED_WIRE_698));


OneBitAdder	b2v_inst341(
	.ci(SYNTHESIZED_WIRE_797),
	.a(SYNTHESIZED_WIRE_798),
	.b(SYNTHESIZED_WIRE_799),
	.co(SYNTHESIZED_WIRE_800),
	.s(SYNTHESIZED_WIRE_701));


OneBitAdder	b2v_inst342(
	.ci(SYNTHESIZED_WIRE_800),
	.a(SYNTHESIZED_WIRE_801),
	.b(SYNTHESIZED_WIRE_802),
	.co(SYNTHESIZED_WIRE_803),
	.s(SYNTHESIZED_WIRE_704));


OneBitAdder	b2v_inst343(
	.ci(SYNTHESIZED_WIRE_803),
	.a(SYNTHESIZED_WIRE_804),
	.b(SYNTHESIZED_WIRE_805),
	.co(SYNTHESIZED_WIRE_806),
	.s(SYNTHESIZED_WIRE_707));


OneBitAdder	b2v_inst344(
	.ci(SYNTHESIZED_WIRE_806),
	.a(SYNTHESIZED_WIRE_807),
	.b(SYNTHESIZED_WIRE_808),
	.co(SYNTHESIZED_WIRE_809),
	.s(SYNTHESIZED_WIRE_710));


OneBitAdder	b2v_inst345(
	.ci(SYNTHESIZED_WIRE_809),
	.a(SYNTHESIZED_WIRE_810),
	.b(SYNTHESIZED_WIRE_811),
	.co(SYNTHESIZED_WIRE_812),
	.s(SYNTHESIZED_WIRE_713));


OneBitAdder	b2v_inst346(
	.ci(SYNTHESIZED_WIRE_812),
	.a(SYNTHESIZED_WIRE_813),
	.b(SYNTHESIZED_WIRE_814),
	.co(SYNTHESIZED_WIRE_815),
	.s(SYNTHESIZED_WIRE_716));


OneBitAdder	b2v_inst347(
	.ci(SYNTHESIZED_WIRE_815),
	.a(SYNTHESIZED_WIRE_816),
	.b(SYNTHESIZED_WIRE_817),
	.co(SYNTHESIZED_WIRE_818),
	.s(SYNTHESIZED_WIRE_719));


OneBitAdder	b2v_inst348(
	.ci(SYNTHESIZED_WIRE_818),
	.a(SYNTHESIZED_WIRE_819),
	.b(SYNTHESIZED_WIRE_820),
	.co(SYNTHESIZED_WIRE_821),
	.s(SYNTHESIZED_WIRE_722));


OneBitAdder	b2v_inst349(
	.ci(SYNTHESIZED_WIRE_821),
	.a(SYNTHESIZED_WIRE_822),
	.b(SYNTHESIZED_WIRE_823),
	.co(SYNTHESIZED_WIRE_827),
	.s(SYNTHESIZED_WIRE_725));


OneBitAdder	b2v_inst35(
	.ci(SYNTHESIZED_WIRE_824),
	.a(SYNTHESIZED_WIRE_825),
	.b(SYNTHESIZED_WIRE_826),
	.co(SYNTHESIZED_WIRE_856),
	.s(Z_ALTERA_SYNTHESIZED[48]));


OneBitAdder	b2v_inst350(
	.ci(SYNTHESIZED_WIRE_827),
	.a(SYNTHESIZED_WIRE_828),
	.b(SYNTHESIZED_WIRE_829),
	.co(SYNTHESIZED_WIRE_830),
	.s(SYNTHESIZED_WIRE_728));


OneBitAdder	b2v_inst351(
	.ci(SYNTHESIZED_WIRE_830),
	.a(SYNTHESIZED_WIRE_831),
	.b(SYNTHESIZED_WIRE_832),
	.co(SYNTHESIZED_WIRE_833),
	.s(SYNTHESIZED_WIRE_731));


OneBitAdder	b2v_inst352(
	.ci(SYNTHESIZED_WIRE_833),
	.a(SYNTHESIZED_WIRE_834),
	.b(SYNTHESIZED_WIRE_835),
	.co(SYNTHESIZED_WIRE_740),
	.s(SYNTHESIZED_WIRE_734));


OneBitAdderHalf	b2v_inst353(
	.A(SYNTHESIZED_WIRE_836),
	.B(SYNTHESIZED_WIRE_837),
	.C(SYNTHESIZED_WIRE_886),
	.S(Z_ALTERA_SYNTHESIZED[21]));


OneBitAdder	b2v_inst354(
	.ci(SYNTHESIZED_WIRE_838),
	.a(SYNTHESIZED_WIRE_839),
	.b(SYNTHESIZED_WIRE_840),
	.co(SYNTHESIZED_WIRE_841),
	.s(SYNTHESIZED_WIRE_835));


OneBitAdder	b2v_inst355(
	.ci(SYNTHESIZED_WIRE_841),
	.a(SYNTHESIZED_WIRE_842),
	.b(SYNTHESIZED_WIRE_843),
	.co(SYNTHESIZED_WIRE_844),
	.s(SYNTHESIZED_WIRE_742));


OneBitAdder	b2v_inst356(
	.ci(SYNTHESIZED_WIRE_844),
	.a(SYNTHESIZED_WIRE_845),
	.b(SYNTHESIZED_WIRE_846),
	.co(SYNTHESIZED_WIRE_847),
	.s(SYNTHESIZED_WIRE_745));


OneBitAdder	b2v_inst357(
	.ci(SYNTHESIZED_WIRE_847),
	.a(SYNTHESIZED_WIRE_848),
	.b(SYNTHESIZED_WIRE_849),
	.co(SYNTHESIZED_WIRE_850),
	.s(SYNTHESIZED_WIRE_748));


OneBitAdder	b2v_inst358(
	.ci(SYNTHESIZED_WIRE_850),
	.a(SYNTHESIZED_WIRE_851),
	.b(SYNTHESIZED_WIRE_852),
	.co(SYNTHESIZED_WIRE_853),
	.s(SYNTHESIZED_WIRE_751));


OneBitAdder	b2v_inst359(
	.ci(SYNTHESIZED_WIRE_853),
	.a(SYNTHESIZED_WIRE_854),
	.b(SYNTHESIZED_WIRE_855),
	.co(SYNTHESIZED_WIRE_859),
	.s(SYNTHESIZED_WIRE_754));


OneBitAdder	b2v_inst36(
	.ci(SYNTHESIZED_WIRE_856),
	.a(SYNTHESIZED_WIRE_857),
	.b(SYNTHESIZED_WIRE_858),
	.co(SYNTHESIZED_WIRE_889),
	.s(Z_ALTERA_SYNTHESIZED[49]));


OneBitAdder	b2v_inst360(
	.ci(SYNTHESIZED_WIRE_859),
	.a(SYNTHESIZED_WIRE_860),
	.b(SYNTHESIZED_WIRE_861),
	.co(SYNTHESIZED_WIRE_862),
	.s(SYNTHESIZED_WIRE_757));


OneBitAdder	b2v_inst361(
	.ci(SYNTHESIZED_WIRE_862),
	.a(SYNTHESIZED_WIRE_863),
	.b(SYNTHESIZED_WIRE_864),
	.co(SYNTHESIZED_WIRE_865),
	.s(SYNTHESIZED_WIRE_760));


OneBitAdder	b2v_inst362(
	.ci(SYNTHESIZED_WIRE_865),
	.a(SYNTHESIZED_WIRE_866),
	.b(SYNTHESIZED_WIRE_867),
	.co(SYNTHESIZED_WIRE_868),
	.s(SYNTHESIZED_WIRE_763));


OneBitAdder	b2v_inst363(
	.ci(SYNTHESIZED_WIRE_868),
	.a(SYNTHESIZED_WIRE_869),
	.b(SYNTHESIZED_WIRE_870),
	.co(SYNTHESIZED_WIRE_871),
	.s(SYNTHESIZED_WIRE_766));


OneBitAdder	b2v_inst364(
	.ci(SYNTHESIZED_WIRE_871),
	.a(SYNTHESIZED_WIRE_872),
	.b(SYNTHESIZED_WIRE_873),
	.co(SYNTHESIZED_WIRE_874),
	.s(SYNTHESIZED_WIRE_769));


OneBitAdder	b2v_inst365(
	.ci(SYNTHESIZED_WIRE_874),
	.a(SYNTHESIZED_WIRE_875),
	.b(SYNTHESIZED_WIRE_876),
	.co(SYNTHESIZED_WIRE_877),
	.s(SYNTHESIZED_WIRE_772));


OneBitAdder	b2v_inst366(
	.ci(SYNTHESIZED_WIRE_877),
	.a(SYNTHESIZED_WIRE_878),
	.b(SYNTHESIZED_WIRE_879),
	.co(SYNTHESIZED_WIRE_880),
	.s(SYNTHESIZED_WIRE_775));


OneBitAdder	b2v_inst367(
	.ci(SYNTHESIZED_WIRE_880),
	.a(SYNTHESIZED_WIRE_881),
	.b(SYNTHESIZED_WIRE_882),
	.co(SYNTHESIZED_WIRE_883),
	.s(SYNTHESIZED_WIRE_778));


OneBitAdder	b2v_inst368(
	.ci(SYNTHESIZED_WIRE_883),
	.a(SYNTHESIZED_WIRE_884),
	.b(SYNTHESIZED_WIRE_885),
	.co(SYNTHESIZED_WIRE_784),
	.s(SYNTHESIZED_WIRE_781));


OneBitAdder	b2v_inst369(
	.ci(SYNTHESIZED_WIRE_886),
	.a(SYNTHESIZED_WIRE_887),
	.b(SYNTHESIZED_WIRE_888),
	.co(SYNTHESIZED_WIRE_892),
	.s(SYNTHESIZED_WIRE_738));


OneBitAdder	b2v_inst37(
	.ci(SYNTHESIZED_WIRE_889),
	.a(SYNTHESIZED_WIRE_890),
	.b(SYNTHESIZED_WIRE_891),
	.co(SYNTHESIZED_WIRE_922),
	.s(Z_ALTERA_SYNTHESIZED[50]));


OneBitAdder	b2v_inst370(
	.ci(SYNTHESIZED_WIRE_892),
	.a(SYNTHESIZED_WIRE_893),
	.b(SYNTHESIZED_WIRE_894),
	.co(SYNTHESIZED_WIRE_895),
	.s(SYNTHESIZED_WIRE_787));


OneBitAdder	b2v_inst371(
	.ci(SYNTHESIZED_WIRE_895),
	.a(SYNTHESIZED_WIRE_896),
	.b(SYNTHESIZED_WIRE_897),
	.co(SYNTHESIZED_WIRE_898),
	.s(SYNTHESIZED_WIRE_790));


OneBitAdder	b2v_inst372(
	.ci(SYNTHESIZED_WIRE_898),
	.a(SYNTHESIZED_WIRE_899),
	.b(SYNTHESIZED_WIRE_900),
	.co(SYNTHESIZED_WIRE_901),
	.s(SYNTHESIZED_WIRE_793));


OneBitAdder	b2v_inst373(
	.ci(SYNTHESIZED_WIRE_901),
	.a(SYNTHESIZED_WIRE_902),
	.b(SYNTHESIZED_WIRE_903),
	.co(SYNTHESIZED_WIRE_904),
	.s(SYNTHESIZED_WIRE_796));


OneBitAdder	b2v_inst374(
	.ci(SYNTHESIZED_WIRE_904),
	.a(SYNTHESIZED_WIRE_905),
	.b(SYNTHESIZED_WIRE_906),
	.co(SYNTHESIZED_WIRE_907),
	.s(SYNTHESIZED_WIRE_799));


OneBitAdder	b2v_inst375(
	.ci(SYNTHESIZED_WIRE_907),
	.a(SYNTHESIZED_WIRE_908),
	.b(SYNTHESIZED_WIRE_909),
	.co(SYNTHESIZED_WIRE_910),
	.s(SYNTHESIZED_WIRE_802));


OneBitAdder	b2v_inst376(
	.ci(SYNTHESIZED_WIRE_910),
	.a(SYNTHESIZED_WIRE_911),
	.b(SYNTHESIZED_WIRE_912),
	.co(SYNTHESIZED_WIRE_913),
	.s(SYNTHESIZED_WIRE_805));


OneBitAdder	b2v_inst377(
	.ci(SYNTHESIZED_WIRE_913),
	.a(SYNTHESIZED_WIRE_914),
	.b(SYNTHESIZED_WIRE_915),
	.co(SYNTHESIZED_WIRE_916),
	.s(SYNTHESIZED_WIRE_808));


OneBitAdder	b2v_inst378(
	.ci(SYNTHESIZED_WIRE_916),
	.a(SYNTHESIZED_WIRE_917),
	.b(SYNTHESIZED_WIRE_918),
	.co(SYNTHESIZED_WIRE_919),
	.s(SYNTHESIZED_WIRE_811));


OneBitAdder	b2v_inst379(
	.ci(SYNTHESIZED_WIRE_919),
	.a(SYNTHESIZED_WIRE_920),
	.b(SYNTHESIZED_WIRE_921),
	.co(SYNTHESIZED_WIRE_925),
	.s(SYNTHESIZED_WIRE_814));


OneBitAdder	b2v_inst38(
	.ci(SYNTHESIZED_WIRE_922),
	.a(SYNTHESIZED_WIRE_923),
	.b(SYNTHESIZED_WIRE_924),
	.co(SYNTHESIZED_WIRE_954),
	.s(Z_ALTERA_SYNTHESIZED[51]));


OneBitAdder	b2v_inst380(
	.ci(SYNTHESIZED_WIRE_925),
	.a(SYNTHESIZED_WIRE_926),
	.b(SYNTHESIZED_WIRE_927),
	.co(SYNTHESIZED_WIRE_928),
	.s(SYNTHESIZED_WIRE_817));


OneBitAdder	b2v_inst381(
	.ci(SYNTHESIZED_WIRE_928),
	.a(SYNTHESIZED_WIRE_929),
	.b(SYNTHESIZED_WIRE_930),
	.co(SYNTHESIZED_WIRE_931),
	.s(SYNTHESIZED_WIRE_820));


OneBitAdder	b2v_inst382(
	.ci(SYNTHESIZED_WIRE_931),
	.a(SYNTHESIZED_WIRE_932),
	.b(SYNTHESIZED_WIRE_933),
	.co(SYNTHESIZED_WIRE_934),
	.s(SYNTHESIZED_WIRE_823));


OneBitAdder	b2v_inst383(
	.ci(SYNTHESIZED_WIRE_934),
	.a(SYNTHESIZED_WIRE_935),
	.b(SYNTHESIZED_WIRE_936),
	.co(SYNTHESIZED_WIRE_937),
	.s(SYNTHESIZED_WIRE_829));


OneBitAdder	b2v_inst384(
	.ci(SYNTHESIZED_WIRE_937),
	.a(SYNTHESIZED_WIRE_938),
	.b(SYNTHESIZED_WIRE_939),
	.co(SYNTHESIZED_WIRE_838),
	.s(SYNTHESIZED_WIRE_832));


OneBitAdderHalf	b2v_inst385(
	.A(SYNTHESIZED_WIRE_940),
	.B(SYNTHESIZED_WIRE_941),
	.C(SYNTHESIZED_WIRE_993),
	.S(Z_ALTERA_SYNTHESIZED[20]));


OneBitAdder	b2v_inst386(
	.ci(SYNTHESIZED_WIRE_942),
	.a(SYNTHESIZED_WIRE_943),
	.b(SYNTHESIZED_WIRE_944),
	.co(SYNTHESIZED_WIRE_945),
	.s(SYNTHESIZED_WIRE_939));


OneBitAdder	b2v_inst387(
	.ci(SYNTHESIZED_WIRE_945),
	.a(SYNTHESIZED_WIRE_946),
	.b(SYNTHESIZED_WIRE_947),
	.co(SYNTHESIZED_WIRE_948),
	.s(SYNTHESIZED_WIRE_840));


OneBitAdder	b2v_inst388(
	.ci(SYNTHESIZED_WIRE_948),
	.a(SYNTHESIZED_WIRE_949),
	.b(SYNTHESIZED_WIRE_950),
	.co(SYNTHESIZED_WIRE_951),
	.s(SYNTHESIZED_WIRE_843));


OneBitAdder	b2v_inst389(
	.ci(SYNTHESIZED_WIRE_951),
	.a(SYNTHESIZED_WIRE_952),
	.b(SYNTHESIZED_WIRE_953),
	.co(SYNTHESIZED_WIRE_957),
	.s(SYNTHESIZED_WIRE_846));


OneBitAdder	b2v_inst39(
	.ci(SYNTHESIZED_WIRE_954),
	.a(SYNTHESIZED_WIRE_955),
	.b(SYNTHESIZED_WIRE_956),
	.co(SYNTHESIZED_WIRE_987),
	.s(Z_ALTERA_SYNTHESIZED[52]));


OneBitAdder	b2v_inst390(
	.ci(SYNTHESIZED_WIRE_957),
	.a(SYNTHESIZED_WIRE_958),
	.b(SYNTHESIZED_WIRE_959),
	.co(SYNTHESIZED_WIRE_960),
	.s(SYNTHESIZED_WIRE_849));


OneBitAdder	b2v_inst391(
	.ci(SYNTHESIZED_WIRE_960),
	.a(SYNTHESIZED_WIRE_961),
	.b(SYNTHESIZED_WIRE_962),
	.co(SYNTHESIZED_WIRE_963),
	.s(SYNTHESIZED_WIRE_852));


OneBitAdder	b2v_inst392(
	.ci(SYNTHESIZED_WIRE_963),
	.a(SYNTHESIZED_WIRE_964),
	.b(SYNTHESIZED_WIRE_965),
	.co(SYNTHESIZED_WIRE_966),
	.s(SYNTHESIZED_WIRE_855));


OneBitAdder	b2v_inst393(
	.ci(SYNTHESIZED_WIRE_966),
	.a(SYNTHESIZED_WIRE_967),
	.b(SYNTHESIZED_WIRE_968),
	.co(SYNTHESIZED_WIRE_969),
	.s(SYNTHESIZED_WIRE_861));


OneBitAdder	b2v_inst394(
	.ci(SYNTHESIZED_WIRE_969),
	.a(SYNTHESIZED_WIRE_970),
	.b(SYNTHESIZED_WIRE_971),
	.co(SYNTHESIZED_WIRE_972),
	.s(SYNTHESIZED_WIRE_864));


OneBitAdder	b2v_inst395(
	.ci(SYNTHESIZED_WIRE_972),
	.a(SYNTHESIZED_WIRE_973),
	.b(SYNTHESIZED_WIRE_974),
	.co(SYNTHESIZED_WIRE_975),
	.s(SYNTHESIZED_WIRE_867));


OneBitAdder	b2v_inst396(
	.ci(SYNTHESIZED_WIRE_975),
	.a(SYNTHESIZED_WIRE_976),
	.b(SYNTHESIZED_WIRE_977),
	.co(SYNTHESIZED_WIRE_978),
	.s(SYNTHESIZED_WIRE_870));


OneBitAdder	b2v_inst397(
	.ci(SYNTHESIZED_WIRE_978),
	.a(SYNTHESIZED_WIRE_979),
	.b(SYNTHESIZED_WIRE_980),
	.co(SYNTHESIZED_WIRE_981),
	.s(SYNTHESIZED_WIRE_873));


OneBitAdder	b2v_inst398(
	.ci(SYNTHESIZED_WIRE_981),
	.a(SYNTHESIZED_WIRE_982),
	.b(SYNTHESIZED_WIRE_983),
	.co(SYNTHESIZED_WIRE_984),
	.s(SYNTHESIZED_WIRE_876));


OneBitAdder	b2v_inst399(
	.ci(SYNTHESIZED_WIRE_984),
	.a(SYNTHESIZED_WIRE_985),
	.b(SYNTHESIZED_WIRE_986),
	.co(SYNTHESIZED_WIRE_990),
	.s(SYNTHESIZED_WIRE_879));


OneBitAdder	b2v_inst40(
	.ci(SYNTHESIZED_WIRE_987),
	.a(SYNTHESIZED_WIRE_988),
	.b(SYNTHESIZED_WIRE_989),
	.co(SYNTHESIZED_WIRE_1020),
	.s(Z_ALTERA_SYNTHESIZED[53]));


OneBitAdder	b2v_inst400(
	.ci(SYNTHESIZED_WIRE_990),
	.a(SYNTHESIZED_WIRE_991),
	.b(SYNTHESIZED_WIRE_992),
	.co(SYNTHESIZED_WIRE_885),
	.s(SYNTHESIZED_WIRE_882));


OneBitAdder	b2v_inst401(
	.ci(SYNTHESIZED_WIRE_993),
	.a(SYNTHESIZED_WIRE_994),
	.b(SYNTHESIZED_WIRE_995),
	.co(SYNTHESIZED_WIRE_996),
	.s(SYNTHESIZED_WIRE_836));


OneBitAdder	b2v_inst402(
	.ci(SYNTHESIZED_WIRE_996),
	.a(SYNTHESIZED_WIRE_997),
	.b(SYNTHESIZED_WIRE_998),
	.co(SYNTHESIZED_WIRE_999),
	.s(SYNTHESIZED_WIRE_888));


OneBitAdder	b2v_inst403(
	.ci(SYNTHESIZED_WIRE_999),
	.a(SYNTHESIZED_WIRE_1000),
	.b(SYNTHESIZED_WIRE_1001),
	.co(SYNTHESIZED_WIRE_1002),
	.s(SYNTHESIZED_WIRE_894));


OneBitAdder	b2v_inst404(
	.ci(SYNTHESIZED_WIRE_1002),
	.a(SYNTHESIZED_WIRE_1003),
	.b(SYNTHESIZED_WIRE_1004),
	.co(SYNTHESIZED_WIRE_1005),
	.s(SYNTHESIZED_WIRE_897));


OneBitAdder	b2v_inst405(
	.ci(SYNTHESIZED_WIRE_1005),
	.a(SYNTHESIZED_WIRE_1006),
	.b(SYNTHESIZED_WIRE_1007),
	.co(SYNTHESIZED_WIRE_1008),
	.s(SYNTHESIZED_WIRE_900));


OneBitAdder	b2v_inst406(
	.ci(SYNTHESIZED_WIRE_1008),
	.a(SYNTHESIZED_WIRE_1009),
	.b(SYNTHESIZED_WIRE_1010),
	.co(SYNTHESIZED_WIRE_1011),
	.s(SYNTHESIZED_WIRE_903));


OneBitAdder	b2v_inst407(
	.ci(SYNTHESIZED_WIRE_1011),
	.a(SYNTHESIZED_WIRE_1012),
	.b(SYNTHESIZED_WIRE_1013),
	.co(SYNTHESIZED_WIRE_1014),
	.s(SYNTHESIZED_WIRE_906));


OneBitAdder	b2v_inst408(
	.ci(SYNTHESIZED_WIRE_1014),
	.a(SYNTHESIZED_WIRE_1015),
	.b(SYNTHESIZED_WIRE_1016),
	.co(SYNTHESIZED_WIRE_1017),
	.s(SYNTHESIZED_WIRE_909));


OneBitAdder	b2v_inst409(
	.ci(SYNTHESIZED_WIRE_1017),
	.a(SYNTHESIZED_WIRE_1018),
	.b(SYNTHESIZED_WIRE_1019),
	.co(SYNTHESIZED_WIRE_1023),
	.s(SYNTHESIZED_WIRE_912));


OneBitAdder	b2v_inst41(
	.ci(SYNTHESIZED_WIRE_1020),
	.a(SYNTHESIZED_WIRE_1021),
	.b(SYNTHESIZED_WIRE_1022),
	.co(SYNTHESIZED_WIRE_1052),
	.s(Z_ALTERA_SYNTHESIZED[54]));


OneBitAdder	b2v_inst410(
	.ci(SYNTHESIZED_WIRE_1023),
	.a(SYNTHESIZED_WIRE_1024),
	.b(SYNTHESIZED_WIRE_1025),
	.co(SYNTHESIZED_WIRE_1026),
	.s(SYNTHESIZED_WIRE_915));


OneBitAdder	b2v_inst411(
	.ci(SYNTHESIZED_WIRE_1026),
	.a(SYNTHESIZED_WIRE_1027),
	.b(SYNTHESIZED_WIRE_1028),
	.co(SYNTHESIZED_WIRE_1029),
	.s(SYNTHESIZED_WIRE_918));


OneBitAdder	b2v_inst412(
	.ci(SYNTHESIZED_WIRE_1029),
	.a(SYNTHESIZED_WIRE_1030),
	.b(SYNTHESIZED_WIRE_1031),
	.co(SYNTHESIZED_WIRE_1032),
	.s(SYNTHESIZED_WIRE_921));


OneBitAdder	b2v_inst413(
	.ci(SYNTHESIZED_WIRE_1032),
	.a(SYNTHESIZED_WIRE_1033),
	.b(SYNTHESIZED_WIRE_1034),
	.co(SYNTHESIZED_WIRE_1035),
	.s(SYNTHESIZED_WIRE_927));


OneBitAdder	b2v_inst414(
	.ci(SYNTHESIZED_WIRE_1035),
	.a(SYNTHESIZED_WIRE_1036),
	.b(SYNTHESIZED_WIRE_1037),
	.co(SYNTHESIZED_WIRE_1038),
	.s(SYNTHESIZED_WIRE_930));


OneBitAdder	b2v_inst415(
	.ci(SYNTHESIZED_WIRE_1038),
	.a(SYNTHESIZED_WIRE_1039),
	.b(SYNTHESIZED_WIRE_1040),
	.co(SYNTHESIZED_WIRE_1041),
	.s(SYNTHESIZED_WIRE_933));


OneBitAdder	b2v_inst416(
	.ci(SYNTHESIZED_WIRE_1041),
	.a(SYNTHESIZED_WIRE_1042),
	.b(SYNTHESIZED_WIRE_1043),
	.co(SYNTHESIZED_WIRE_942),
	.s(SYNTHESIZED_WIRE_936));


OneBitAdderHalf	b2v_inst417(
	.A(SYNTHESIZED_WIRE_1044),
	.B(SYNTHESIZED_WIRE_1045),
	.C(SYNTHESIZED_WIRE_1097),
	.S(Z_ALTERA_SYNTHESIZED[19]));


OneBitAdder	b2v_inst418(
	.ci(SYNTHESIZED_WIRE_1046),
	.a(SYNTHESIZED_WIRE_1047),
	.b(SYNTHESIZED_WIRE_1048),
	.co(SYNTHESIZED_WIRE_1049),
	.s(SYNTHESIZED_WIRE_1043));


OneBitAdder	b2v_inst419(
	.ci(SYNTHESIZED_WIRE_1049),
	.a(SYNTHESIZED_WIRE_1050),
	.b(SYNTHESIZED_WIRE_1051),
	.co(SYNTHESIZED_WIRE_1055),
	.s(SYNTHESIZED_WIRE_944));


OneBitAdder	b2v_inst42(
	.ci(SYNTHESIZED_WIRE_1052),
	.a(SYNTHESIZED_WIRE_1053),
	.b(SYNTHESIZED_WIRE_1054),
	.co(SYNTHESIZED_WIRE_1085),
	.s(Z_ALTERA_SYNTHESIZED[55]));


OneBitAdder	b2v_inst420(
	.ci(SYNTHESIZED_WIRE_1055),
	.a(SYNTHESIZED_WIRE_1056),
	.b(SYNTHESIZED_WIRE_1057),
	.co(SYNTHESIZED_WIRE_1058),
	.s(SYNTHESIZED_WIRE_947));


OneBitAdder	b2v_inst421(
	.ci(SYNTHESIZED_WIRE_1058),
	.a(SYNTHESIZED_WIRE_1059),
	.b(SYNTHESIZED_WIRE_1060),
	.co(SYNTHESIZED_WIRE_1061),
	.s(SYNTHESIZED_WIRE_950));


OneBitAdder	b2v_inst422(
	.ci(SYNTHESIZED_WIRE_1061),
	.a(SYNTHESIZED_WIRE_1062),
	.b(SYNTHESIZED_WIRE_1063),
	.co(SYNTHESIZED_WIRE_1064),
	.s(SYNTHESIZED_WIRE_953));


OneBitAdder	b2v_inst423(
	.ci(SYNTHESIZED_WIRE_1064),
	.a(SYNTHESIZED_WIRE_1065),
	.b(SYNTHESIZED_WIRE_1066),
	.co(SYNTHESIZED_WIRE_1067),
	.s(SYNTHESIZED_WIRE_959));


OneBitAdder	b2v_inst424(
	.ci(SYNTHESIZED_WIRE_1067),
	.a(SYNTHESIZED_WIRE_1068),
	.b(SYNTHESIZED_WIRE_1069),
	.co(SYNTHESIZED_WIRE_1070),
	.s(SYNTHESIZED_WIRE_962));


OneBitAdder	b2v_inst425(
	.ci(SYNTHESIZED_WIRE_1070),
	.a(SYNTHESIZED_WIRE_1071),
	.b(SYNTHESIZED_WIRE_1072),
	.co(SYNTHESIZED_WIRE_1073),
	.s(SYNTHESIZED_WIRE_965));


OneBitAdder	b2v_inst426(
	.ci(SYNTHESIZED_WIRE_1073),
	.a(SYNTHESIZED_WIRE_1074),
	.b(SYNTHESIZED_WIRE_1075),
	.co(SYNTHESIZED_WIRE_1076),
	.s(SYNTHESIZED_WIRE_968));


OneBitAdder	b2v_inst427(
	.ci(SYNTHESIZED_WIRE_1076),
	.a(SYNTHESIZED_WIRE_1077),
	.b(SYNTHESIZED_WIRE_1078),
	.co(SYNTHESIZED_WIRE_1079),
	.s(SYNTHESIZED_WIRE_971));


OneBitAdder	b2v_inst428(
	.ci(SYNTHESIZED_WIRE_1079),
	.a(SYNTHESIZED_WIRE_1080),
	.b(SYNTHESIZED_WIRE_1081),
	.co(SYNTHESIZED_WIRE_1082),
	.s(SYNTHESIZED_WIRE_974));


OneBitAdder	b2v_inst429(
	.ci(SYNTHESIZED_WIRE_1082),
	.a(SYNTHESIZED_WIRE_1083),
	.b(SYNTHESIZED_WIRE_1084),
	.co(SYNTHESIZED_WIRE_1088),
	.s(SYNTHESIZED_WIRE_977));


OneBitAdder	b2v_inst43(
	.ci(SYNTHESIZED_WIRE_1085),
	.a(SYNTHESIZED_WIRE_1086),
	.b(SYNTHESIZED_WIRE_1087),
	.co(SYNTHESIZED_WIRE_1118),
	.s(Z_ALTERA_SYNTHESIZED[56]));


OneBitAdder	b2v_inst430(
	.ci(SYNTHESIZED_WIRE_1088),
	.a(SYNTHESIZED_WIRE_1089),
	.b(SYNTHESIZED_WIRE_1090),
	.co(SYNTHESIZED_WIRE_1091),
	.s(SYNTHESIZED_WIRE_980));


OneBitAdder	b2v_inst431(
	.ci(SYNTHESIZED_WIRE_1091),
	.a(SYNTHESIZED_WIRE_1092),
	.b(SYNTHESIZED_WIRE_1093),
	.co(SYNTHESIZED_WIRE_1094),
	.s(SYNTHESIZED_WIRE_983));


OneBitAdder	b2v_inst432(
	.ci(SYNTHESIZED_WIRE_1094),
	.a(SYNTHESIZED_WIRE_1095),
	.b(SYNTHESIZED_WIRE_1096),
	.co(SYNTHESIZED_WIRE_992),
	.s(SYNTHESIZED_WIRE_986));


OneBitAdder	b2v_inst433(
	.ci(SYNTHESIZED_WIRE_1097),
	.a(SYNTHESIZED_WIRE_1098),
	.b(SYNTHESIZED_WIRE_1099),
	.co(SYNTHESIZED_WIRE_1100),
	.s(SYNTHESIZED_WIRE_940));


OneBitAdder	b2v_inst434(
	.ci(SYNTHESIZED_WIRE_1100),
	.a(SYNTHESIZED_WIRE_1101),
	.b(SYNTHESIZED_WIRE_1102),
	.co(SYNTHESIZED_WIRE_1103),
	.s(SYNTHESIZED_WIRE_995));


OneBitAdder	b2v_inst435(
	.ci(SYNTHESIZED_WIRE_1103),
	.a(SYNTHESIZED_WIRE_1104),
	.b(SYNTHESIZED_WIRE_1105),
	.co(SYNTHESIZED_WIRE_1106),
	.s(SYNTHESIZED_WIRE_998));


OneBitAdder	b2v_inst436(
	.ci(SYNTHESIZED_WIRE_1106),
	.a(SYNTHESIZED_WIRE_1107),
	.b(SYNTHESIZED_WIRE_1108),
	.co(SYNTHESIZED_WIRE_1109),
	.s(SYNTHESIZED_WIRE_1001));


OneBitAdder	b2v_inst437(
	.ci(SYNTHESIZED_WIRE_1109),
	.a(SYNTHESIZED_WIRE_1110),
	.b(SYNTHESIZED_WIRE_1111),
	.co(SYNTHESIZED_WIRE_1112),
	.s(SYNTHESIZED_WIRE_1004));


OneBitAdder	b2v_inst438(
	.ci(SYNTHESIZED_WIRE_1112),
	.a(SYNTHESIZED_WIRE_1113),
	.b(SYNTHESIZED_WIRE_1114),
	.co(SYNTHESIZED_WIRE_1115),
	.s(SYNTHESIZED_WIRE_1007));


OneBitAdder	b2v_inst439(
	.ci(SYNTHESIZED_WIRE_1115),
	.a(SYNTHESIZED_WIRE_1116),
	.b(SYNTHESIZED_WIRE_1117),
	.co(SYNTHESIZED_WIRE_1121),
	.s(SYNTHESIZED_WIRE_1010));


OneBitAdder	b2v_inst44(
	.ci(SYNTHESIZED_WIRE_1118),
	.a(SYNTHESIZED_WIRE_1119),
	.b(SYNTHESIZED_WIRE_1120),
	.co(SYNTHESIZED_WIRE_1150),
	.s(Z_ALTERA_SYNTHESIZED[57]));


OneBitAdder	b2v_inst440(
	.ci(SYNTHESIZED_WIRE_1121),
	.a(SYNTHESIZED_WIRE_1122),
	.b(SYNTHESIZED_WIRE_1123),
	.co(SYNTHESIZED_WIRE_1124),
	.s(SYNTHESIZED_WIRE_1013));


OneBitAdder	b2v_inst441(
	.ci(SYNTHESIZED_WIRE_1124),
	.a(SYNTHESIZED_WIRE_1125),
	.b(SYNTHESIZED_WIRE_1126),
	.co(SYNTHESIZED_WIRE_1127),
	.s(SYNTHESIZED_WIRE_1016));


OneBitAdder	b2v_inst442(
	.ci(SYNTHESIZED_WIRE_1127),
	.a(SYNTHESIZED_WIRE_1128),
	.b(SYNTHESIZED_WIRE_1129),
	.co(SYNTHESIZED_WIRE_1130),
	.s(SYNTHESIZED_WIRE_1019));


OneBitAdder	b2v_inst443(
	.ci(SYNTHESIZED_WIRE_1130),
	.a(SYNTHESIZED_WIRE_1131),
	.b(SYNTHESIZED_WIRE_1132),
	.co(SYNTHESIZED_WIRE_1133),
	.s(SYNTHESIZED_WIRE_1025));


OneBitAdder	b2v_inst444(
	.ci(SYNTHESIZED_WIRE_1133),
	.a(SYNTHESIZED_WIRE_1134),
	.b(SYNTHESIZED_WIRE_1135),
	.co(SYNTHESIZED_WIRE_1136),
	.s(SYNTHESIZED_WIRE_1028));


OneBitAdder	b2v_inst445(
	.ci(SYNTHESIZED_WIRE_1136),
	.a(SYNTHESIZED_WIRE_1137),
	.b(SYNTHESIZED_WIRE_1138),
	.co(SYNTHESIZED_WIRE_1139),
	.s(SYNTHESIZED_WIRE_1031));


OneBitAdder	b2v_inst446(
	.ci(SYNTHESIZED_WIRE_1139),
	.a(SYNTHESIZED_WIRE_1140),
	.b(SYNTHESIZED_WIRE_1141),
	.co(SYNTHESIZED_WIRE_1142),
	.s(SYNTHESIZED_WIRE_1034));


OneBitAdder	b2v_inst447(
	.ci(SYNTHESIZED_WIRE_1142),
	.a(SYNTHESIZED_WIRE_1143),
	.b(SYNTHESIZED_WIRE_1144),
	.co(SYNTHESIZED_WIRE_1145),
	.s(SYNTHESIZED_WIRE_1037));


OneBitAdder	b2v_inst448(
	.ci(SYNTHESIZED_WIRE_1145),
	.a(SYNTHESIZED_WIRE_1146),
	.b(SYNTHESIZED_WIRE_1147),
	.co(SYNTHESIZED_WIRE_1046),
	.s(SYNTHESIZED_WIRE_1040));


OneBitAdderHalf	b2v_inst449(
	.A(SYNTHESIZED_WIRE_1148),
	.B(SYNTHESIZED_WIRE_1149),
	.C(SYNTHESIZED_WIRE_1201),
	.S(Z_ALTERA_SYNTHESIZED[18]));


OneBitAdder	b2v_inst45(
	.ci(SYNTHESIZED_WIRE_1150),
	.a(SYNTHESIZED_WIRE_1151),
	.b(SYNTHESIZED_WIRE_1152),
	.co(SYNTHESIZED_WIRE_1183),
	.s(Z_ALTERA_SYNTHESIZED[58]));


OneBitAdder	b2v_inst450(
	.ci(SYNTHESIZED_WIRE_1153),
	.a(SYNTHESIZED_WIRE_1154),
	.b(SYNTHESIZED_WIRE_1155),
	.co(SYNTHESIZED_WIRE_1156),
	.s(SYNTHESIZED_WIRE_1147));


OneBitAdder	b2v_inst451(
	.ci(SYNTHESIZED_WIRE_1156),
	.a(SYNTHESIZED_WIRE_1157),
	.b(SYNTHESIZED_WIRE_1158),
	.co(SYNTHESIZED_WIRE_1159),
	.s(SYNTHESIZED_WIRE_1048));


OneBitAdder	b2v_inst452(
	.ci(SYNTHESIZED_WIRE_1159),
	.a(SYNTHESIZED_WIRE_1160),
	.b(SYNTHESIZED_WIRE_1161),
	.co(SYNTHESIZED_WIRE_1162),
	.s(SYNTHESIZED_WIRE_1051));


OneBitAdder	b2v_inst453(
	.ci(SYNTHESIZED_WIRE_1162),
	.a(SYNTHESIZED_WIRE_1163),
	.b(SYNTHESIZED_WIRE_1164),
	.co(SYNTHESIZED_WIRE_1165),
	.s(SYNTHESIZED_WIRE_1057));


OneBitAdder	b2v_inst454(
	.ci(SYNTHESIZED_WIRE_1165),
	.a(SYNTHESIZED_WIRE_1166),
	.b(SYNTHESIZED_WIRE_1167),
	.co(SYNTHESIZED_WIRE_1168),
	.s(SYNTHESIZED_WIRE_1060));


OneBitAdder	b2v_inst455(
	.ci(SYNTHESIZED_WIRE_1168),
	.a(SYNTHESIZED_WIRE_1169),
	.b(SYNTHESIZED_WIRE_1170),
	.co(SYNTHESIZED_WIRE_1171),
	.s(SYNTHESIZED_WIRE_1063));


OneBitAdder	b2v_inst456(
	.ci(SYNTHESIZED_WIRE_1171),
	.a(SYNTHESIZED_WIRE_1172),
	.b(SYNTHESIZED_WIRE_1173),
	.co(SYNTHESIZED_WIRE_1174),
	.s(SYNTHESIZED_WIRE_1066));


OneBitAdder	b2v_inst457(
	.ci(SYNTHESIZED_WIRE_1174),
	.a(SYNTHESIZED_WIRE_1175),
	.b(SYNTHESIZED_WIRE_1176),
	.co(SYNTHESIZED_WIRE_1177),
	.s(SYNTHESIZED_WIRE_1069));


OneBitAdder	b2v_inst458(
	.ci(SYNTHESIZED_WIRE_1177),
	.a(SYNTHESIZED_WIRE_1178),
	.b(SYNTHESIZED_WIRE_1179),
	.co(SYNTHESIZED_WIRE_1180),
	.s(SYNTHESIZED_WIRE_1072));


OneBitAdder	b2v_inst459(
	.ci(SYNTHESIZED_WIRE_1180),
	.a(SYNTHESIZED_WIRE_1181),
	.b(SYNTHESIZED_WIRE_1182),
	.co(SYNTHESIZED_WIRE_1186),
	.s(SYNTHESIZED_WIRE_1075));


OneBitAdder	b2v_inst46(
	.ci(SYNTHESIZED_WIRE_1183),
	.a(SYNTHESIZED_WIRE_1184),
	.b(SYNTHESIZED_WIRE_1185),
	.co(SYNTHESIZED_WIRE_1216),
	.s(Z_ALTERA_SYNTHESIZED[59]));


OneBitAdder	b2v_inst460(
	.ci(SYNTHESIZED_WIRE_1186),
	.a(SYNTHESIZED_WIRE_1187),
	.b(SYNTHESIZED_WIRE_1188),
	.co(SYNTHESIZED_WIRE_1189),
	.s(SYNTHESIZED_WIRE_1078));


OneBitAdder	b2v_inst461(
	.ci(SYNTHESIZED_WIRE_1189),
	.a(SYNTHESIZED_WIRE_1190),
	.b(SYNTHESIZED_WIRE_1191),
	.co(SYNTHESIZED_WIRE_1192),
	.s(SYNTHESIZED_WIRE_1081));


OneBitAdder	b2v_inst462(
	.ci(SYNTHESIZED_WIRE_1192),
	.a(SYNTHESIZED_WIRE_1193),
	.b(SYNTHESIZED_WIRE_1194),
	.co(SYNTHESIZED_WIRE_1195),
	.s(SYNTHESIZED_WIRE_1084));


OneBitAdder	b2v_inst463(
	.ci(SYNTHESIZED_WIRE_1195),
	.a(SYNTHESIZED_WIRE_1196),
	.b(SYNTHESIZED_WIRE_1197),
	.co(SYNTHESIZED_WIRE_1198),
	.s(SYNTHESIZED_WIRE_1090));


OneBitAdder	b2v_inst464(
	.ci(SYNTHESIZED_WIRE_1198),
	.a(SYNTHESIZED_WIRE_1199),
	.b(SYNTHESIZED_WIRE_1200),
	.co(SYNTHESIZED_WIRE_1096),
	.s(SYNTHESIZED_WIRE_1093));


OneBitAdder	b2v_inst465(
	.ci(SYNTHESIZED_WIRE_1201),
	.a(SYNTHESIZED_WIRE_1202),
	.b(SYNTHESIZED_WIRE_1203),
	.co(SYNTHESIZED_WIRE_1204),
	.s(SYNTHESIZED_WIRE_1044));


OneBitAdder	b2v_inst466(
	.ci(SYNTHESIZED_WIRE_1204),
	.a(SYNTHESIZED_WIRE_1205),
	.b(SYNTHESIZED_WIRE_1206),
	.co(SYNTHESIZED_WIRE_1207),
	.s(SYNTHESIZED_WIRE_1099));


OneBitAdder	b2v_inst467(
	.ci(SYNTHESIZED_WIRE_1207),
	.a(SYNTHESIZED_WIRE_1208),
	.b(SYNTHESIZED_WIRE_1209),
	.co(SYNTHESIZED_WIRE_1210),
	.s(SYNTHESIZED_WIRE_1102));


OneBitAdder	b2v_inst468(
	.ci(SYNTHESIZED_WIRE_1210),
	.a(SYNTHESIZED_WIRE_1211),
	.b(SYNTHESIZED_WIRE_1212),
	.co(SYNTHESIZED_WIRE_1213),
	.s(SYNTHESIZED_WIRE_1105));


OneBitAdder	b2v_inst469(
	.ci(SYNTHESIZED_WIRE_1213),
	.a(SYNTHESIZED_WIRE_1214),
	.b(SYNTHESIZED_WIRE_1215),
	.co(SYNTHESIZED_WIRE_1219),
	.s(SYNTHESIZED_WIRE_1108));


OneBitAdder	b2v_inst47(
	.ci(SYNTHESIZED_WIRE_1216),
	.a(SYNTHESIZED_WIRE_1217),
	.b(SYNTHESIZED_WIRE_1218),
	.co(SYNTHESIZED_WIRE_1249),
	.s(Z_ALTERA_SYNTHESIZED[60]));


OneBitAdder	b2v_inst470(
	.ci(SYNTHESIZED_WIRE_1219),
	.a(SYNTHESIZED_WIRE_1220),
	.b(SYNTHESIZED_WIRE_1221),
	.co(SYNTHESIZED_WIRE_1222),
	.s(SYNTHESIZED_WIRE_1111));


OneBitAdder	b2v_inst471(
	.ci(SYNTHESIZED_WIRE_1222),
	.a(SYNTHESIZED_WIRE_1223),
	.b(SYNTHESIZED_WIRE_1224),
	.co(SYNTHESIZED_WIRE_1225),
	.s(SYNTHESIZED_WIRE_1114));


OneBitAdder	b2v_inst472(
	.ci(SYNTHESIZED_WIRE_1225),
	.a(SYNTHESIZED_WIRE_1226),
	.b(SYNTHESIZED_WIRE_1227),
	.co(SYNTHESIZED_WIRE_1228),
	.s(SYNTHESIZED_WIRE_1117));


OneBitAdder	b2v_inst473(
	.ci(SYNTHESIZED_WIRE_1228),
	.a(SYNTHESIZED_WIRE_1229),
	.b(SYNTHESIZED_WIRE_1230),
	.co(SYNTHESIZED_WIRE_1231),
	.s(SYNTHESIZED_WIRE_1123));


OneBitAdder	b2v_inst474(
	.ci(SYNTHESIZED_WIRE_1231),
	.a(SYNTHESIZED_WIRE_1232),
	.b(SYNTHESIZED_WIRE_1233),
	.co(SYNTHESIZED_WIRE_1234),
	.s(SYNTHESIZED_WIRE_1126));


OneBitAdder	b2v_inst475(
	.ci(SYNTHESIZED_WIRE_1234),
	.a(SYNTHESIZED_WIRE_1235),
	.b(SYNTHESIZED_WIRE_1236),
	.co(SYNTHESIZED_WIRE_1237),
	.s(SYNTHESIZED_WIRE_1129));


OneBitAdder	b2v_inst476(
	.ci(SYNTHESIZED_WIRE_1237),
	.a(SYNTHESIZED_WIRE_1238),
	.b(SYNTHESIZED_WIRE_1239),
	.co(SYNTHESIZED_WIRE_1240),
	.s(SYNTHESIZED_WIRE_1132));


OneBitAdder	b2v_inst477(
	.ci(SYNTHESIZED_WIRE_1240),
	.a(SYNTHESIZED_WIRE_1241),
	.b(SYNTHESIZED_WIRE_1242),
	.co(SYNTHESIZED_WIRE_1243),
	.s(SYNTHESIZED_WIRE_1135));


OneBitAdder	b2v_inst478(
	.ci(SYNTHESIZED_WIRE_1243),
	.a(SYNTHESIZED_WIRE_1244),
	.b(SYNTHESIZED_WIRE_1245),
	.co(SYNTHESIZED_WIRE_1246),
	.s(SYNTHESIZED_WIRE_1138));


OneBitAdder	b2v_inst479(
	.ci(SYNTHESIZED_WIRE_1246),
	.a(SYNTHESIZED_WIRE_1247),
	.b(SYNTHESIZED_WIRE_1248),
	.co(SYNTHESIZED_WIRE_1252),
	.s(SYNTHESIZED_WIRE_1141));


OneBitAdder	b2v_inst48(
	.ci(SYNTHESIZED_WIRE_1249),
	.a(SYNTHESIZED_WIRE_1250),
	.b(SYNTHESIZED_WIRE_1251),
	.co(SYNTHESIZED_WIRE_1281),
	.s(Z_ALTERA_SYNTHESIZED[61]));


OneBitAdder	b2v_inst480(
	.ci(SYNTHESIZED_WIRE_1252),
	.a(SYNTHESIZED_WIRE_1253),
	.b(SYNTHESIZED_WIRE_1254),
	.co(SYNTHESIZED_WIRE_1153),
	.s(SYNTHESIZED_WIRE_1144));


OneBitAdderHalf	b2v_inst481(
	.A(SYNTHESIZED_WIRE_1255),
	.B(SYNTHESIZED_WIRE_1256),
	.C(SYNTHESIZED_WIRE_1305),
	.S(Z_ALTERA_SYNTHESIZED[17]));


OneBitAdder	b2v_inst482(
	.ci(SYNTHESIZED_WIRE_1257),
	.a(SYNTHESIZED_WIRE_1258),
	.b(SYNTHESIZED_WIRE_1259),
	.co(SYNTHESIZED_WIRE_1260),
	.s(SYNTHESIZED_WIRE_1254));


OneBitAdder	b2v_inst483(
	.ci(SYNTHESIZED_WIRE_1260),
	.a(SYNTHESIZED_WIRE_1261),
	.b(SYNTHESIZED_WIRE_1262),
	.co(SYNTHESIZED_WIRE_1263),
	.s(SYNTHESIZED_WIRE_1155));


OneBitAdder	b2v_inst484(
	.ci(SYNTHESIZED_WIRE_1263),
	.a(SYNTHESIZED_WIRE_1264),
	.b(SYNTHESIZED_WIRE_1265),
	.co(SYNTHESIZED_WIRE_1266),
	.s(SYNTHESIZED_WIRE_1158));


OneBitAdder	b2v_inst485(
	.ci(SYNTHESIZED_WIRE_1266),
	.a(SYNTHESIZED_WIRE_1267),
	.b(SYNTHESIZED_WIRE_1268),
	.co(SYNTHESIZED_WIRE_1269),
	.s(SYNTHESIZED_WIRE_1161));


OneBitAdder	b2v_inst486(
	.ci(SYNTHESIZED_WIRE_1269),
	.a(SYNTHESIZED_WIRE_1270),
	.b(SYNTHESIZED_WIRE_1271),
	.co(SYNTHESIZED_WIRE_1272),
	.s(SYNTHESIZED_WIRE_1164));


OneBitAdder	b2v_inst487(
	.ci(SYNTHESIZED_WIRE_1272),
	.a(SYNTHESIZED_WIRE_1273),
	.b(SYNTHESIZED_WIRE_1274),
	.co(SYNTHESIZED_WIRE_1275),
	.s(SYNTHESIZED_WIRE_1167));


OneBitAdder	b2v_inst488(
	.ci(SYNTHESIZED_WIRE_1275),
	.a(SYNTHESIZED_WIRE_1276),
	.b(SYNTHESIZED_WIRE_1277),
	.co(SYNTHESIZED_WIRE_1278),
	.s(SYNTHESIZED_WIRE_1170));


OneBitAdder	b2v_inst489(
	.ci(SYNTHESIZED_WIRE_1278),
	.a(SYNTHESIZED_WIRE_1279),
	.b(SYNTHESIZED_WIRE_1280),
	.co(SYNTHESIZED_WIRE_1284),
	.s(SYNTHESIZED_WIRE_1173));


OneBitAdder	b2v_inst49(
	.ci(SYNTHESIZED_WIRE_1281),
	.a(SYNTHESIZED_WIRE_1282),
	.b(SYNTHESIZED_WIRE_1283),
	.co(SYNTHESIZED_WIRE_673),
	.s(Z_ALTERA_SYNTHESIZED[62]));


OneBitAdder	b2v_inst490(
	.ci(SYNTHESIZED_WIRE_1284),
	.a(SYNTHESIZED_WIRE_1285),
	.b(SYNTHESIZED_WIRE_1286),
	.co(SYNTHESIZED_WIRE_1287),
	.s(SYNTHESIZED_WIRE_1176));


OneBitAdder	b2v_inst491(
	.ci(SYNTHESIZED_WIRE_1287),
	.a(SYNTHESIZED_WIRE_1288),
	.b(SYNTHESIZED_WIRE_1289),
	.co(SYNTHESIZED_WIRE_1290),
	.s(SYNTHESIZED_WIRE_1179));


OneBitAdder	b2v_inst492(
	.ci(SYNTHESIZED_WIRE_1290),
	.a(SYNTHESIZED_WIRE_1291),
	.b(SYNTHESIZED_WIRE_1292),
	.co(SYNTHESIZED_WIRE_1293),
	.s(SYNTHESIZED_WIRE_1182));


OneBitAdder	b2v_inst493(
	.ci(SYNTHESIZED_WIRE_1293),
	.a(SYNTHESIZED_WIRE_1294),
	.b(SYNTHESIZED_WIRE_1295),
	.co(SYNTHESIZED_WIRE_1296),
	.s(SYNTHESIZED_WIRE_1188));


OneBitAdder	b2v_inst494(
	.ci(SYNTHESIZED_WIRE_1296),
	.a(SYNTHESIZED_WIRE_1297),
	.b(SYNTHESIZED_WIRE_1298),
	.co(SYNTHESIZED_WIRE_1299),
	.s(SYNTHESIZED_WIRE_1191));


OneBitAdder	b2v_inst495(
	.ci(SYNTHESIZED_WIRE_1299),
	.a(SYNTHESIZED_WIRE_1300),
	.b(SYNTHESIZED_WIRE_1301),
	.co(SYNTHESIZED_WIRE_1302),
	.s(SYNTHESIZED_WIRE_1194));


OneBitAdder	b2v_inst496(
	.ci(SYNTHESIZED_WIRE_1302),
	.a(SYNTHESIZED_WIRE_1303),
	.b(SYNTHESIZED_WIRE_1304),
	.co(SYNTHESIZED_WIRE_1200),
	.s(SYNTHESIZED_WIRE_1197));


OneBitAdder	b2v_inst497(
	.ci(SYNTHESIZED_WIRE_1305),
	.a(SYNTHESIZED_WIRE_1306),
	.b(SYNTHESIZED_WIRE_1307),
	.co(SYNTHESIZED_WIRE_1308),
	.s(SYNTHESIZED_WIRE_1148));


OneBitAdder	b2v_inst498(
	.ci(SYNTHESIZED_WIRE_1308),
	.a(SYNTHESIZED_WIRE_1309),
	.b(SYNTHESIZED_WIRE_1310),
	.co(SYNTHESIZED_WIRE_1311),
	.s(SYNTHESIZED_WIRE_1203));


OneBitAdder	b2v_inst499(
	.ci(SYNTHESIZED_WIRE_1311),
	.a(SYNTHESIZED_WIRE_1312),
	.b(SYNTHESIZED_WIRE_1313),
	.co(SYNTHESIZED_WIRE_1317),
	.s(SYNTHESIZED_WIRE_1206));


OneBitAdder	b2v_inst50(
	.ci(SYNTHESIZED_WIRE_1314),
	.a(SYNTHESIZED_WIRE_1315),
	.b(SYNTHESIZED_WIRE_1316),
	.co(SYNTHESIZED_WIRE_1347),
	.s(Z_ALTERA_SYNTHESIZED[32]));


OneBitAdder	b2v_inst500(
	.ci(SYNTHESIZED_WIRE_1317),
	.a(SYNTHESIZED_WIRE_1318),
	.b(SYNTHESIZED_WIRE_1319),
	.co(SYNTHESIZED_WIRE_1320),
	.s(SYNTHESIZED_WIRE_1209));


OneBitAdder	b2v_inst501(
	.ci(SYNTHESIZED_WIRE_1320),
	.a(SYNTHESIZED_WIRE_1321),
	.b(SYNTHESIZED_WIRE_1322),
	.co(SYNTHESIZED_WIRE_1323),
	.s(SYNTHESIZED_WIRE_1212));


OneBitAdder	b2v_inst502(
	.ci(SYNTHESIZED_WIRE_1323),
	.a(SYNTHESIZED_WIRE_1324),
	.b(SYNTHESIZED_WIRE_1325),
	.co(SYNTHESIZED_WIRE_1326),
	.s(SYNTHESIZED_WIRE_1215));


OneBitAdder	b2v_inst503(
	.ci(SYNTHESIZED_WIRE_1326),
	.a(SYNTHESIZED_WIRE_1327),
	.b(SYNTHESIZED_WIRE_1328),
	.co(SYNTHESIZED_WIRE_1329),
	.s(SYNTHESIZED_WIRE_1221));


OneBitAdder	b2v_inst504(
	.ci(SYNTHESIZED_WIRE_1329),
	.a(SYNTHESIZED_WIRE_1330),
	.b(SYNTHESIZED_WIRE_1331),
	.co(SYNTHESIZED_WIRE_1332),
	.s(SYNTHESIZED_WIRE_1224));


OneBitAdder	b2v_inst505(
	.ci(SYNTHESIZED_WIRE_1332),
	.a(SYNTHESIZED_WIRE_1333),
	.b(SYNTHESIZED_WIRE_1334),
	.co(SYNTHESIZED_WIRE_1335),
	.s(SYNTHESIZED_WIRE_1227));


OneBitAdder	b2v_inst506(
	.ci(SYNTHESIZED_WIRE_1335),
	.a(SYNTHESIZED_WIRE_1336),
	.b(SYNTHESIZED_WIRE_1337),
	.co(SYNTHESIZED_WIRE_1338),
	.s(SYNTHESIZED_WIRE_1230));


OneBitAdder	b2v_inst507(
	.ci(SYNTHESIZED_WIRE_1338),
	.a(SYNTHESIZED_WIRE_1339),
	.b(SYNTHESIZED_WIRE_1340),
	.co(SYNTHESIZED_WIRE_1341),
	.s(SYNTHESIZED_WIRE_1233));


OneBitAdder	b2v_inst508(
	.ci(SYNTHESIZED_WIRE_1341),
	.a(SYNTHESIZED_WIRE_1342),
	.b(SYNTHESIZED_WIRE_1343),
	.co(SYNTHESIZED_WIRE_1344),
	.s(SYNTHESIZED_WIRE_1236));


OneBitAdder	b2v_inst509(
	.ci(SYNTHESIZED_WIRE_1344),
	.a(SYNTHESIZED_WIRE_1345),
	.b(SYNTHESIZED_WIRE_1346),
	.co(SYNTHESIZED_WIRE_1350),
	.s(SYNTHESIZED_WIRE_1239));


OneBitAdder	b2v_inst51(
	.ci(SYNTHESIZED_WIRE_1347),
	.a(SYNTHESIZED_WIRE_1348),
	.b(SYNTHESIZED_WIRE_1349),
	.co(SYNTHESIZED_WIRE_1379),
	.s(Z_ALTERA_SYNTHESIZED[33]));


OneBitAdder	b2v_inst510(
	.ci(SYNTHESIZED_WIRE_1350),
	.a(SYNTHESIZED_WIRE_1351),
	.b(SYNTHESIZED_WIRE_1352),
	.co(SYNTHESIZED_WIRE_1353),
	.s(SYNTHESIZED_WIRE_1242));


OneBitAdder	b2v_inst511(
	.ci(SYNTHESIZED_WIRE_1353),
	.a(SYNTHESIZED_WIRE_1354),
	.b(SYNTHESIZED_WIRE_1355),
	.co(SYNTHESIZED_WIRE_1356),
	.s(SYNTHESIZED_WIRE_1245));


OneBitAdder	b2v_inst512(
	.ci(SYNTHESIZED_WIRE_1356),
	.a(SYNTHESIZED_WIRE_1357),
	.b(SYNTHESIZED_WIRE_1358),
	.co(SYNTHESIZED_WIRE_1257),
	.s(SYNTHESIZED_WIRE_1248));


OneBitAdderHalf	b2v_inst513(
	.A(SYNTHESIZED_WIRE_1359),
	.B(SYNTHESIZED_WIRE_1360),
	.C(SYNTHESIZED_WIRE_1409),
	.S(Z_ALTERA_SYNTHESIZED[16]));


OneBitAdder	b2v_inst514(
	.ci(SYNTHESIZED_WIRE_1361),
	.a(SYNTHESIZED_WIRE_1362),
	.b(SYNTHESIZED_WIRE_1363),
	.co(SYNTHESIZED_WIRE_1364),
	.s(SYNTHESIZED_WIRE_1358));


OneBitAdder	b2v_inst515(
	.ci(SYNTHESIZED_WIRE_1364),
	.a(SYNTHESIZED_WIRE_1365),
	.b(SYNTHESIZED_WIRE_1366),
	.co(SYNTHESIZED_WIRE_1367),
	.s(SYNTHESIZED_WIRE_1259));


OneBitAdder	b2v_inst516(
	.ci(SYNTHESIZED_WIRE_1367),
	.a(SYNTHESIZED_WIRE_1368),
	.b(SYNTHESIZED_WIRE_1369),
	.co(SYNTHESIZED_WIRE_1370),
	.s(SYNTHESIZED_WIRE_1262));


OneBitAdder	b2v_inst517(
	.ci(SYNTHESIZED_WIRE_1370),
	.a(SYNTHESIZED_WIRE_1371),
	.b(SYNTHESIZED_WIRE_1372),
	.co(SYNTHESIZED_WIRE_1373),
	.s(SYNTHESIZED_WIRE_1265));


OneBitAdder	b2v_inst518(
	.ci(SYNTHESIZED_WIRE_1373),
	.a(SYNTHESIZED_WIRE_1374),
	.b(SYNTHESIZED_WIRE_1375),
	.co(SYNTHESIZED_WIRE_1376),
	.s(SYNTHESIZED_WIRE_1268));


OneBitAdder	b2v_inst519(
	.ci(SYNTHESIZED_WIRE_1376),
	.a(SYNTHESIZED_WIRE_1377),
	.b(SYNTHESIZED_WIRE_1378),
	.co(SYNTHESIZED_WIRE_1382),
	.s(SYNTHESIZED_WIRE_1271));


OneBitAdder	b2v_inst52(
	.ci(SYNTHESIZED_WIRE_1379),
	.a(SYNTHESIZED_WIRE_1380),
	.b(SYNTHESIZED_WIRE_1381),
	.co(SYNTHESIZED_WIRE_1412),
	.s(Z_ALTERA_SYNTHESIZED[34]));


OneBitAdder	b2v_inst520(
	.ci(SYNTHESIZED_WIRE_1382),
	.a(SYNTHESIZED_WIRE_1383),
	.b(SYNTHESIZED_WIRE_1384),
	.co(SYNTHESIZED_WIRE_1385),
	.s(SYNTHESIZED_WIRE_1274));


OneBitAdder	b2v_inst521(
	.ci(SYNTHESIZED_WIRE_1385),
	.a(SYNTHESIZED_WIRE_1386),
	.b(SYNTHESIZED_WIRE_1387),
	.co(SYNTHESIZED_WIRE_1388),
	.s(SYNTHESIZED_WIRE_1277));


OneBitAdder	b2v_inst522(
	.ci(SYNTHESIZED_WIRE_1388),
	.a(SYNTHESIZED_WIRE_1389),
	.b(SYNTHESIZED_WIRE_1390),
	.co(SYNTHESIZED_WIRE_1391),
	.s(SYNTHESIZED_WIRE_1280));


OneBitAdder	b2v_inst523(
	.ci(SYNTHESIZED_WIRE_1391),
	.a(SYNTHESIZED_WIRE_1392),
	.b(SYNTHESIZED_WIRE_1393),
	.co(SYNTHESIZED_WIRE_1394),
	.s(SYNTHESIZED_WIRE_1286));


OneBitAdder	b2v_inst524(
	.ci(SYNTHESIZED_WIRE_1394),
	.a(SYNTHESIZED_WIRE_1395),
	.b(SYNTHESIZED_WIRE_1396),
	.co(SYNTHESIZED_WIRE_1397),
	.s(SYNTHESIZED_WIRE_1289));


OneBitAdder	b2v_inst525(
	.ci(SYNTHESIZED_WIRE_1397),
	.a(SYNTHESIZED_WIRE_1398),
	.b(SYNTHESIZED_WIRE_1399),
	.co(SYNTHESIZED_WIRE_1400),
	.s(SYNTHESIZED_WIRE_1292));


OneBitAdder	b2v_inst526(
	.ci(SYNTHESIZED_WIRE_1400),
	.a(SYNTHESIZED_WIRE_1401),
	.b(SYNTHESIZED_WIRE_1402),
	.co(SYNTHESIZED_WIRE_1403),
	.s(SYNTHESIZED_WIRE_1295));


OneBitAdder	b2v_inst527(
	.ci(SYNTHESIZED_WIRE_1403),
	.a(SYNTHESIZED_WIRE_1404),
	.b(SYNTHESIZED_WIRE_1405),
	.co(SYNTHESIZED_WIRE_1406),
	.s(SYNTHESIZED_WIRE_1298));


OneBitAdder	b2v_inst528(
	.ci(SYNTHESIZED_WIRE_1406),
	.a(SYNTHESIZED_WIRE_1407),
	.b(SYNTHESIZED_WIRE_1408),
	.co(SYNTHESIZED_WIRE_1304),
	.s(SYNTHESIZED_WIRE_1301));


OneBitAdder	b2v_inst529(
	.ci(SYNTHESIZED_WIRE_1409),
	.a(SYNTHESIZED_WIRE_1410),
	.b(SYNTHESIZED_WIRE_1411),
	.co(SYNTHESIZED_WIRE_1415),
	.s(SYNTHESIZED_WIRE_1255));


OneBitAdder	b2v_inst53(
	.ci(SYNTHESIZED_WIRE_1412),
	.a(SYNTHESIZED_WIRE_1413),
	.b(SYNTHESIZED_WIRE_1414),
	.co(SYNTHESIZED_WIRE_1445),
	.s(Z_ALTERA_SYNTHESIZED[35]));


OneBitAdder	b2v_inst530(
	.ci(SYNTHESIZED_WIRE_1415),
	.a(SYNTHESIZED_WIRE_1416),
	.b(SYNTHESIZED_WIRE_1417),
	.co(SYNTHESIZED_WIRE_1418),
	.s(SYNTHESIZED_WIRE_1307));


OneBitAdder	b2v_inst531(
	.ci(SYNTHESIZED_WIRE_1418),
	.a(SYNTHESIZED_WIRE_1419),
	.b(SYNTHESIZED_WIRE_1420),
	.co(SYNTHESIZED_WIRE_1421),
	.s(SYNTHESIZED_WIRE_1310));


OneBitAdder	b2v_inst532(
	.ci(SYNTHESIZED_WIRE_1421),
	.a(SYNTHESIZED_WIRE_1422),
	.b(SYNTHESIZED_WIRE_1423),
	.co(SYNTHESIZED_WIRE_1424),
	.s(SYNTHESIZED_WIRE_1313));


OneBitAdder	b2v_inst533(
	.ci(SYNTHESIZED_WIRE_1424),
	.a(SYNTHESIZED_WIRE_1425),
	.b(SYNTHESIZED_WIRE_1426),
	.co(SYNTHESIZED_WIRE_1427),
	.s(SYNTHESIZED_WIRE_1319));


OneBitAdder	b2v_inst534(
	.ci(SYNTHESIZED_WIRE_1427),
	.a(SYNTHESIZED_WIRE_1428),
	.b(SYNTHESIZED_WIRE_1429),
	.co(SYNTHESIZED_WIRE_1430),
	.s(SYNTHESIZED_WIRE_1322));


OneBitAdder	b2v_inst535(
	.ci(SYNTHESIZED_WIRE_1430),
	.a(SYNTHESIZED_WIRE_1431),
	.b(SYNTHESIZED_WIRE_1432),
	.co(SYNTHESIZED_WIRE_1433),
	.s(SYNTHESIZED_WIRE_1325));


OneBitAdder	b2v_inst536(
	.ci(SYNTHESIZED_WIRE_1433),
	.a(SYNTHESIZED_WIRE_1434),
	.b(SYNTHESIZED_WIRE_1435),
	.co(SYNTHESIZED_WIRE_1436),
	.s(SYNTHESIZED_WIRE_1328));


OneBitAdder	b2v_inst537(
	.ci(SYNTHESIZED_WIRE_1436),
	.a(SYNTHESIZED_WIRE_1437),
	.b(SYNTHESIZED_WIRE_1438),
	.co(SYNTHESIZED_WIRE_1439),
	.s(SYNTHESIZED_WIRE_1331));


OneBitAdder	b2v_inst538(
	.ci(SYNTHESIZED_WIRE_1439),
	.a(SYNTHESIZED_WIRE_1440),
	.b(SYNTHESIZED_WIRE_1441),
	.co(SYNTHESIZED_WIRE_1442),
	.s(SYNTHESIZED_WIRE_1334));


OneBitAdder	b2v_inst539(
	.ci(SYNTHESIZED_WIRE_1442),
	.a(SYNTHESIZED_WIRE_1443),
	.b(SYNTHESIZED_WIRE_1444),
	.co(SYNTHESIZED_WIRE_1448),
	.s(SYNTHESIZED_WIRE_1337));


OneBitAdder	b2v_inst54(
	.ci(SYNTHESIZED_WIRE_1445),
	.a(SYNTHESIZED_WIRE_1446),
	.b(SYNTHESIZED_WIRE_1447),
	.co(SYNTHESIZED_WIRE_1477),
	.s(Z_ALTERA_SYNTHESIZED[36]));


OneBitAdder	b2v_inst540(
	.ci(SYNTHESIZED_WIRE_1448),
	.a(SYNTHESIZED_WIRE_1449),
	.b(SYNTHESIZED_WIRE_1450),
	.co(SYNTHESIZED_WIRE_1451),
	.s(SYNTHESIZED_WIRE_1340));


OneBitAdder	b2v_inst541(
	.ci(SYNTHESIZED_WIRE_1451),
	.a(SYNTHESIZED_WIRE_1452),
	.b(SYNTHESIZED_WIRE_1453),
	.co(SYNTHESIZED_WIRE_1454),
	.s(SYNTHESIZED_WIRE_1343));


OneBitAdder	b2v_inst542(
	.ci(SYNTHESIZED_WIRE_1454),
	.a(SYNTHESIZED_WIRE_1455),
	.b(SYNTHESIZED_WIRE_1456),
	.co(SYNTHESIZED_WIRE_1457),
	.s(SYNTHESIZED_WIRE_1346));


OneBitAdder	b2v_inst543(
	.ci(SYNTHESIZED_WIRE_1457),
	.a(SYNTHESIZED_WIRE_1458),
	.b(SYNTHESIZED_WIRE_1459),
	.co(SYNTHESIZED_WIRE_1460),
	.s(SYNTHESIZED_WIRE_1352));


OneBitAdder	b2v_inst544(
	.ci(SYNTHESIZED_WIRE_1460),
	.a(SYNTHESIZED_WIRE_1461),
	.b(SYNTHESIZED_WIRE_1462),
	.co(SYNTHESIZED_WIRE_1361),
	.s(SYNTHESIZED_WIRE_1355));


OneBitAdderHalf	b2v_inst545(
	.A(SYNTHESIZED_WIRE_1463),
	.B(SYNTHESIZED_WIRE_1464),
	.C(SYNTHESIZED_WIRE_1516),
	.S(Z_ALTERA_SYNTHESIZED[15]));


OneBitAdder	b2v_inst546(
	.ci(SYNTHESIZED_WIRE_1465),
	.a(SYNTHESIZED_WIRE_1466),
	.b(SYNTHESIZED_WIRE_1467),
	.co(SYNTHESIZED_WIRE_1468),
	.s(SYNTHESIZED_WIRE_1462));


OneBitAdder	b2v_inst547(
	.ci(SYNTHESIZED_WIRE_1468),
	.a(SYNTHESIZED_WIRE_1469),
	.b(SYNTHESIZED_WIRE_1470),
	.co(SYNTHESIZED_WIRE_1471),
	.s(SYNTHESIZED_WIRE_1363));


OneBitAdder	b2v_inst548(
	.ci(SYNTHESIZED_WIRE_1471),
	.a(SYNTHESIZED_WIRE_1472),
	.b(SYNTHESIZED_WIRE_1473),
	.co(SYNTHESIZED_WIRE_1474),
	.s(SYNTHESIZED_WIRE_1366));


OneBitAdder	b2v_inst549(
	.ci(SYNTHESIZED_WIRE_1474),
	.a(SYNTHESIZED_WIRE_1475),
	.b(SYNTHESIZED_WIRE_1476),
	.co(SYNTHESIZED_WIRE_1480),
	.s(SYNTHESIZED_WIRE_1369));


OneBitAdder	b2v_inst55(
	.ci(SYNTHESIZED_WIRE_1477),
	.a(SYNTHESIZED_WIRE_1478),
	.b(SYNTHESIZED_WIRE_1479),
	.co(SYNTHESIZED_WIRE_1510),
	.s(Z_ALTERA_SYNTHESIZED[37]));


OneBitAdder	b2v_inst550(
	.ci(SYNTHESIZED_WIRE_1480),
	.a(SYNTHESIZED_WIRE_1481),
	.b(SYNTHESIZED_WIRE_1482),
	.co(SYNTHESIZED_WIRE_1483),
	.s(SYNTHESIZED_WIRE_1372));


OneBitAdder	b2v_inst551(
	.ci(SYNTHESIZED_WIRE_1483),
	.a(SYNTHESIZED_WIRE_1484),
	.b(SYNTHESIZED_WIRE_1485),
	.co(SYNTHESIZED_WIRE_1486),
	.s(SYNTHESIZED_WIRE_1375));


OneBitAdder	b2v_inst552(
	.ci(SYNTHESIZED_WIRE_1486),
	.a(SYNTHESIZED_WIRE_1487),
	.b(SYNTHESIZED_WIRE_1488),
	.co(SYNTHESIZED_WIRE_1489),
	.s(SYNTHESIZED_WIRE_1378));


OneBitAdder	b2v_inst553(
	.ci(SYNTHESIZED_WIRE_1489),
	.a(SYNTHESIZED_WIRE_1490),
	.b(SYNTHESIZED_WIRE_1491),
	.co(SYNTHESIZED_WIRE_1492),
	.s(SYNTHESIZED_WIRE_1384));


OneBitAdder	b2v_inst554(
	.ci(SYNTHESIZED_WIRE_1492),
	.a(SYNTHESIZED_WIRE_1493),
	.b(SYNTHESIZED_WIRE_1494),
	.co(SYNTHESIZED_WIRE_1495),
	.s(SYNTHESIZED_WIRE_1387));


OneBitAdder	b2v_inst555(
	.ci(SYNTHESIZED_WIRE_1495),
	.a(SYNTHESIZED_WIRE_1496),
	.b(SYNTHESIZED_WIRE_1497),
	.co(SYNTHESIZED_WIRE_1498),
	.s(SYNTHESIZED_WIRE_1390));


OneBitAdder	b2v_inst556(
	.ci(SYNTHESIZED_WIRE_1498),
	.a(SYNTHESIZED_WIRE_1499),
	.b(SYNTHESIZED_WIRE_1500),
	.co(SYNTHESIZED_WIRE_1501),
	.s(SYNTHESIZED_WIRE_1393));


OneBitAdder	b2v_inst557(
	.ci(SYNTHESIZED_WIRE_1501),
	.a(SYNTHESIZED_WIRE_1502),
	.b(SYNTHESIZED_WIRE_1503),
	.co(SYNTHESIZED_WIRE_1504),
	.s(SYNTHESIZED_WIRE_1396));


OneBitAdder	b2v_inst558(
	.ci(SYNTHESIZED_WIRE_1504),
	.a(SYNTHESIZED_WIRE_1505),
	.b(SYNTHESIZED_WIRE_1506),
	.co(SYNTHESIZED_WIRE_1507),
	.s(SYNTHESIZED_WIRE_1399));


OneBitAdder	b2v_inst559(
	.ci(SYNTHESIZED_WIRE_1507),
	.a(SYNTHESIZED_WIRE_1508),
	.b(SYNTHESIZED_WIRE_1509),
	.co(SYNTHESIZED_WIRE_1513),
	.s(SYNTHESIZED_WIRE_1402));


OneBitAdder	b2v_inst56(
	.ci(SYNTHESIZED_WIRE_1510),
	.a(SYNTHESIZED_WIRE_1511),
	.b(SYNTHESIZED_WIRE_1512),
	.co(SYNTHESIZED_WIRE_1543),
	.s(Z_ALTERA_SYNTHESIZED[38]));


OneBitAdder	b2v_inst560(
	.ci(SYNTHESIZED_WIRE_1513),
	.a(SYNTHESIZED_WIRE_1514),
	.b(SYNTHESIZED_WIRE_1515),
	.co(SYNTHESIZED_WIRE_1408),
	.s(SYNTHESIZED_WIRE_1405));


OneBitAdder	b2v_inst561(
	.ci(SYNTHESIZED_WIRE_1516),
	.a(SYNTHESIZED_WIRE_1517),
	.b(SYNTHESIZED_WIRE_1518),
	.co(SYNTHESIZED_WIRE_1519),
	.s(SYNTHESIZED_WIRE_1359));


OneBitAdder	b2v_inst562(
	.ci(SYNTHESIZED_WIRE_1519),
	.a(SYNTHESIZED_WIRE_1520),
	.b(SYNTHESIZED_WIRE_1521),
	.co(SYNTHESIZED_WIRE_1522),
	.s(SYNTHESIZED_WIRE_1411));


OneBitAdder	b2v_inst563(
	.ci(SYNTHESIZED_WIRE_1522),
	.a(SYNTHESIZED_WIRE_1523),
	.b(SYNTHESIZED_WIRE_1524),
	.co(SYNTHESIZED_WIRE_1525),
	.s(SYNTHESIZED_WIRE_1417));


OneBitAdder	b2v_inst564(
	.ci(SYNTHESIZED_WIRE_1525),
	.a(SYNTHESIZED_WIRE_1526),
	.b(SYNTHESIZED_WIRE_1527),
	.co(SYNTHESIZED_WIRE_1528),
	.s(SYNTHESIZED_WIRE_1420));


OneBitAdder	b2v_inst565(
	.ci(SYNTHESIZED_WIRE_1528),
	.a(SYNTHESIZED_WIRE_1529),
	.b(SYNTHESIZED_WIRE_1530),
	.co(SYNTHESIZED_WIRE_1531),
	.s(SYNTHESIZED_WIRE_1423));


OneBitAdder	b2v_inst566(
	.ci(SYNTHESIZED_WIRE_1531),
	.a(SYNTHESIZED_WIRE_1532),
	.b(SYNTHESIZED_WIRE_1533),
	.co(SYNTHESIZED_WIRE_1534),
	.s(SYNTHESIZED_WIRE_1426));


OneBitAdder	b2v_inst567(
	.ci(SYNTHESIZED_WIRE_1534),
	.a(SYNTHESIZED_WIRE_1535),
	.b(SYNTHESIZED_WIRE_1536),
	.co(SYNTHESIZED_WIRE_1537),
	.s(SYNTHESIZED_WIRE_1429));


OneBitAdder	b2v_inst568(
	.ci(SYNTHESIZED_WIRE_1537),
	.a(SYNTHESIZED_WIRE_1538),
	.b(SYNTHESIZED_WIRE_1539),
	.co(SYNTHESIZED_WIRE_1540),
	.s(SYNTHESIZED_WIRE_1432));


OneBitAdder	b2v_inst569(
	.ci(SYNTHESIZED_WIRE_1540),
	.a(SYNTHESIZED_WIRE_1541),
	.b(SYNTHESIZED_WIRE_1542),
	.co(SYNTHESIZED_WIRE_1546),
	.s(SYNTHESIZED_WIRE_1435));


OneBitAdder	b2v_inst57(
	.ci(SYNTHESIZED_WIRE_1543),
	.a(SYNTHESIZED_WIRE_1544),
	.b(SYNTHESIZED_WIRE_1545),
	.co(SYNTHESIZED_WIRE_1575),
	.s(Z_ALTERA_SYNTHESIZED[39]));


OneBitAdder	b2v_inst570(
	.ci(SYNTHESIZED_WIRE_1546),
	.a(SYNTHESIZED_WIRE_1547),
	.b(SYNTHESIZED_WIRE_1548),
	.co(SYNTHESIZED_WIRE_1549),
	.s(SYNTHESIZED_WIRE_1438));


OneBitAdder	b2v_inst571(
	.ci(SYNTHESIZED_WIRE_1549),
	.a(SYNTHESIZED_WIRE_1550),
	.b(SYNTHESIZED_WIRE_1551),
	.co(SYNTHESIZED_WIRE_1552),
	.s(SYNTHESIZED_WIRE_1441));


OneBitAdder	b2v_inst572(
	.ci(SYNTHESIZED_WIRE_1552),
	.a(SYNTHESIZED_WIRE_1553),
	.b(SYNTHESIZED_WIRE_1554),
	.co(SYNTHESIZED_WIRE_1555),
	.s(SYNTHESIZED_WIRE_1444));


OneBitAdder	b2v_inst573(
	.ci(SYNTHESIZED_WIRE_1555),
	.a(SYNTHESIZED_WIRE_1556),
	.b(SYNTHESIZED_WIRE_1557),
	.co(SYNTHESIZED_WIRE_1558),
	.s(SYNTHESIZED_WIRE_1450));


OneBitAdder	b2v_inst574(
	.ci(SYNTHESIZED_WIRE_1558),
	.a(SYNTHESIZED_WIRE_1559),
	.b(SYNTHESIZED_WIRE_1560),
	.co(SYNTHESIZED_WIRE_1561),
	.s(SYNTHESIZED_WIRE_1453));


OneBitAdder	b2v_inst575(
	.ci(SYNTHESIZED_WIRE_1561),
	.a(SYNTHESIZED_WIRE_1562),
	.b(SYNTHESIZED_WIRE_1563),
	.co(SYNTHESIZED_WIRE_1564),
	.s(SYNTHESIZED_WIRE_1456));


OneBitAdder	b2v_inst576(
	.ci(SYNTHESIZED_WIRE_1564),
	.a(SYNTHESIZED_WIRE_1565),
	.b(SYNTHESIZED_WIRE_1566),
	.co(SYNTHESIZED_WIRE_1465),
	.s(SYNTHESIZED_WIRE_1459));


OneBitAdderHalf	b2v_inst577(
	.A(SYNTHESIZED_WIRE_1567),
	.B(SYNTHESIZED_WIRE_1568),
	.C(SYNTHESIZED_WIRE_1620),
	.S(Z_ALTERA_SYNTHESIZED[14]));


OneBitAdder	b2v_inst578(
	.ci(SYNTHESIZED_WIRE_1569),
	.a(SYNTHESIZED_WIRE_1570),
	.b(SYNTHESIZED_WIRE_1571),
	.co(SYNTHESIZED_WIRE_1572),
	.s(SYNTHESIZED_WIRE_1566));


OneBitAdder	b2v_inst579(
	.ci(SYNTHESIZED_WIRE_1572),
	.a(SYNTHESIZED_WIRE_1573),
	.b(SYNTHESIZED_WIRE_1574),
	.co(SYNTHESIZED_WIRE_1578),
	.s(SYNTHESIZED_WIRE_1467));


OneBitAdder	b2v_inst58(
	.ci(SYNTHESIZED_WIRE_1575),
	.a(SYNTHESIZED_WIRE_1576),
	.b(SYNTHESIZED_WIRE_1577),
	.co(SYNTHESIZED_WIRE_1608),
	.s(Z_ALTERA_SYNTHESIZED[40]));


OneBitAdder	b2v_inst580(
	.ci(SYNTHESIZED_WIRE_1578),
	.a(SYNTHESIZED_WIRE_1579),
	.b(SYNTHESIZED_WIRE_1580),
	.co(SYNTHESIZED_WIRE_1581),
	.s(SYNTHESIZED_WIRE_1470));


OneBitAdder	b2v_inst581(
	.ci(SYNTHESIZED_WIRE_1581),
	.a(SYNTHESIZED_WIRE_1582),
	.b(SYNTHESIZED_WIRE_1583),
	.co(SYNTHESIZED_WIRE_1584),
	.s(SYNTHESIZED_WIRE_1473));


OneBitAdder	b2v_inst582(
	.ci(SYNTHESIZED_WIRE_1584),
	.a(SYNTHESIZED_WIRE_1585),
	.b(SYNTHESIZED_WIRE_1586),
	.co(SYNTHESIZED_WIRE_1587),
	.s(SYNTHESIZED_WIRE_1476));


OneBitAdder	b2v_inst583(
	.ci(SYNTHESIZED_WIRE_1587),
	.a(SYNTHESIZED_WIRE_1588),
	.b(SYNTHESIZED_WIRE_1589),
	.co(SYNTHESIZED_WIRE_1590),
	.s(SYNTHESIZED_WIRE_1482));


OneBitAdder	b2v_inst584(
	.ci(SYNTHESIZED_WIRE_1590),
	.a(SYNTHESIZED_WIRE_1591),
	.b(SYNTHESIZED_WIRE_1592),
	.co(SYNTHESIZED_WIRE_1593),
	.s(SYNTHESIZED_WIRE_1485));


OneBitAdder	b2v_inst585(
	.ci(SYNTHESIZED_WIRE_1593),
	.a(SYNTHESIZED_WIRE_1594),
	.b(SYNTHESIZED_WIRE_1595),
	.co(SYNTHESIZED_WIRE_1596),
	.s(SYNTHESIZED_WIRE_1488));


OneBitAdder	b2v_inst586(
	.ci(SYNTHESIZED_WIRE_1596),
	.a(SYNTHESIZED_WIRE_1597),
	.b(SYNTHESIZED_WIRE_1598),
	.co(SYNTHESIZED_WIRE_1599),
	.s(SYNTHESIZED_WIRE_1491));


OneBitAdder	b2v_inst587(
	.ci(SYNTHESIZED_WIRE_1599),
	.a(SYNTHESIZED_WIRE_1600),
	.b(SYNTHESIZED_WIRE_1601),
	.co(SYNTHESIZED_WIRE_1602),
	.s(SYNTHESIZED_WIRE_1494));


OneBitAdder	b2v_inst588(
	.ci(SYNTHESIZED_WIRE_1602),
	.a(SYNTHESIZED_WIRE_1603),
	.b(SYNTHESIZED_WIRE_1604),
	.co(SYNTHESIZED_WIRE_1605),
	.s(SYNTHESIZED_WIRE_1497));


OneBitAdder	b2v_inst589(
	.ci(SYNTHESIZED_WIRE_1605),
	.a(SYNTHESIZED_WIRE_1606),
	.b(SYNTHESIZED_WIRE_1607),
	.co(SYNTHESIZED_WIRE_1611),
	.s(SYNTHESIZED_WIRE_1500));


OneBitAdder	b2v_inst59(
	.ci(SYNTHESIZED_WIRE_1608),
	.a(SYNTHESIZED_WIRE_1609),
	.b(SYNTHESIZED_WIRE_1610),
	.co(SYNTHESIZED_WIRE_1641),
	.s(Z_ALTERA_SYNTHESIZED[41]));


OneBitAdder	b2v_inst590(
	.ci(SYNTHESIZED_WIRE_1611),
	.a(SYNTHESIZED_WIRE_1612),
	.b(SYNTHESIZED_WIRE_1613),
	.co(SYNTHESIZED_WIRE_1614),
	.s(SYNTHESIZED_WIRE_1503));


OneBitAdder	b2v_inst591(
	.ci(SYNTHESIZED_WIRE_1614),
	.a(SYNTHESIZED_WIRE_1615),
	.b(SYNTHESIZED_WIRE_1616),
	.co(SYNTHESIZED_WIRE_1617),
	.s(SYNTHESIZED_WIRE_1506));


OneBitAdder	b2v_inst592(
	.ci(SYNTHESIZED_WIRE_1617),
	.a(SYNTHESIZED_WIRE_1618),
	.b(SYNTHESIZED_WIRE_1619),
	.co(SYNTHESIZED_WIRE_1515),
	.s(SYNTHESIZED_WIRE_1509));


OneBitAdder	b2v_inst593(
	.ci(SYNTHESIZED_WIRE_1620),
	.a(SYNTHESIZED_WIRE_1621),
	.b(SYNTHESIZED_WIRE_1622),
	.co(SYNTHESIZED_WIRE_1623),
	.s(SYNTHESIZED_WIRE_1463));


OneBitAdder	b2v_inst594(
	.ci(SYNTHESIZED_WIRE_1623),
	.a(SYNTHESIZED_WIRE_1624),
	.b(SYNTHESIZED_WIRE_1625),
	.co(SYNTHESIZED_WIRE_1626),
	.s(SYNTHESIZED_WIRE_1518));


OneBitAdder	b2v_inst595(
	.ci(SYNTHESIZED_WIRE_1626),
	.a(SYNTHESIZED_WIRE_1627),
	.b(SYNTHESIZED_WIRE_1628),
	.co(SYNTHESIZED_WIRE_1629),
	.s(SYNTHESIZED_WIRE_1521));


OneBitAdder	b2v_inst596(
	.ci(SYNTHESIZED_WIRE_1629),
	.a(SYNTHESIZED_WIRE_1630),
	.b(SYNTHESIZED_WIRE_1631),
	.co(SYNTHESIZED_WIRE_1632),
	.s(SYNTHESIZED_WIRE_1524));


OneBitAdder	b2v_inst597(
	.ci(SYNTHESIZED_WIRE_1632),
	.a(SYNTHESIZED_WIRE_1633),
	.b(SYNTHESIZED_WIRE_1634),
	.co(SYNTHESIZED_WIRE_1635),
	.s(SYNTHESIZED_WIRE_1527));


OneBitAdder	b2v_inst598(
	.ci(SYNTHESIZED_WIRE_1635),
	.a(SYNTHESIZED_WIRE_1636),
	.b(SYNTHESIZED_WIRE_1637),
	.co(SYNTHESIZED_WIRE_1638),
	.s(SYNTHESIZED_WIRE_1530));


OneBitAdder	b2v_inst599(
	.ci(SYNTHESIZED_WIRE_1638),
	.a(SYNTHESIZED_WIRE_1639),
	.b(SYNTHESIZED_WIRE_1640),
	.co(SYNTHESIZED_WIRE_1644),
	.s(SYNTHESIZED_WIRE_1533));


OneBitAdder	b2v_inst60(
	.ci(SYNTHESIZED_WIRE_1641),
	.a(SYNTHESIZED_WIRE_1642),
	.b(SYNTHESIZED_WIRE_1643),
	.co(SYNTHESIZED_WIRE_1673),
	.s(Z_ALTERA_SYNTHESIZED[42]));


OneBitAdder	b2v_inst600(
	.ci(SYNTHESIZED_WIRE_1644),
	.a(SYNTHESIZED_WIRE_1645),
	.b(SYNTHESIZED_WIRE_1646),
	.co(SYNTHESIZED_WIRE_1647),
	.s(SYNTHESIZED_WIRE_1536));


OneBitAdder	b2v_inst601(
	.ci(SYNTHESIZED_WIRE_1647),
	.a(SYNTHESIZED_WIRE_1648),
	.b(SYNTHESIZED_WIRE_1649),
	.co(SYNTHESIZED_WIRE_1650),
	.s(SYNTHESIZED_WIRE_1539));


OneBitAdder	b2v_inst602(
	.ci(SYNTHESIZED_WIRE_1650),
	.a(SYNTHESIZED_WIRE_1651),
	.b(SYNTHESIZED_WIRE_1652),
	.co(SYNTHESIZED_WIRE_1653),
	.s(SYNTHESIZED_WIRE_1542));


OneBitAdder	b2v_inst603(
	.ci(SYNTHESIZED_WIRE_1653),
	.a(SYNTHESIZED_WIRE_1654),
	.b(SYNTHESIZED_WIRE_1655),
	.co(SYNTHESIZED_WIRE_1656),
	.s(SYNTHESIZED_WIRE_1548));


OneBitAdder	b2v_inst604(
	.ci(SYNTHESIZED_WIRE_1656),
	.a(SYNTHESIZED_WIRE_1657),
	.b(SYNTHESIZED_WIRE_1658),
	.co(SYNTHESIZED_WIRE_1659),
	.s(SYNTHESIZED_WIRE_1551));


OneBitAdder	b2v_inst605(
	.ci(SYNTHESIZED_WIRE_1659),
	.a(SYNTHESIZED_WIRE_1660),
	.b(SYNTHESIZED_WIRE_1661),
	.co(SYNTHESIZED_WIRE_1662),
	.s(SYNTHESIZED_WIRE_1554));


OneBitAdder	b2v_inst606(
	.ci(SYNTHESIZED_WIRE_1662),
	.a(SYNTHESIZED_WIRE_1663),
	.b(SYNTHESIZED_WIRE_1664),
	.co(SYNTHESIZED_WIRE_1665),
	.s(SYNTHESIZED_WIRE_1557));


OneBitAdder	b2v_inst607(
	.ci(SYNTHESIZED_WIRE_1665),
	.a(SYNTHESIZED_WIRE_1666),
	.b(SYNTHESIZED_WIRE_1667),
	.co(SYNTHESIZED_WIRE_1668),
	.s(SYNTHESIZED_WIRE_1560));


OneBitAdder	b2v_inst608(
	.ci(SYNTHESIZED_WIRE_1668),
	.a(SYNTHESIZED_WIRE_1669),
	.b(SYNTHESIZED_WIRE_1670),
	.co(SYNTHESIZED_WIRE_1569),
	.s(SYNTHESIZED_WIRE_1563));


OneBitAdderHalf	b2v_inst609(
	.A(SYNTHESIZED_WIRE_1671),
	.B(SYNTHESIZED_WIRE_1672),
	.C(SYNTHESIZED_WIRE_1724),
	.S(Z_ALTERA_SYNTHESIZED[13]));


OneBitAdder	b2v_inst61(
	.ci(SYNTHESIZED_WIRE_1673),
	.a(SYNTHESIZED_WIRE_1674),
	.b(SYNTHESIZED_WIRE_1675),
	.co(SYNTHESIZED_WIRE_1706),
	.s(Z_ALTERA_SYNTHESIZED[43]));


OneBitAdder	b2v_inst610(
	.ci(SYNTHESIZED_WIRE_1676),
	.a(SYNTHESIZED_WIRE_1677),
	.b(SYNTHESIZED_WIRE_1678),
	.co(SYNTHESIZED_WIRE_1679),
	.s(SYNTHESIZED_WIRE_1670));


OneBitAdder	b2v_inst611(
	.ci(SYNTHESIZED_WIRE_1679),
	.a(SYNTHESIZED_WIRE_1680),
	.b(SYNTHESIZED_WIRE_1681),
	.co(SYNTHESIZED_WIRE_1682),
	.s(SYNTHESIZED_WIRE_1571));


OneBitAdder	b2v_inst612(
	.ci(SYNTHESIZED_WIRE_1682),
	.a(SYNTHESIZED_WIRE_1683),
	.b(SYNTHESIZED_WIRE_1684),
	.co(SYNTHESIZED_WIRE_1685),
	.s(SYNTHESIZED_WIRE_1574));


OneBitAdder	b2v_inst613(
	.ci(SYNTHESIZED_WIRE_1685),
	.a(SYNTHESIZED_WIRE_1686),
	.b(SYNTHESIZED_WIRE_1687),
	.co(SYNTHESIZED_WIRE_1688),
	.s(SYNTHESIZED_WIRE_1580));


OneBitAdder	b2v_inst614(
	.ci(SYNTHESIZED_WIRE_1688),
	.a(SYNTHESIZED_WIRE_1689),
	.b(SYNTHESIZED_WIRE_1690),
	.co(SYNTHESIZED_WIRE_1691),
	.s(SYNTHESIZED_WIRE_1583));


OneBitAdder	b2v_inst615(
	.ci(SYNTHESIZED_WIRE_1691),
	.a(SYNTHESIZED_WIRE_1692),
	.b(SYNTHESIZED_WIRE_1693),
	.co(SYNTHESIZED_WIRE_1694),
	.s(SYNTHESIZED_WIRE_1586));


OneBitAdder	b2v_inst616(
	.ci(SYNTHESIZED_WIRE_1694),
	.a(SYNTHESIZED_WIRE_1695),
	.b(SYNTHESIZED_WIRE_1696),
	.co(SYNTHESIZED_WIRE_1697),
	.s(SYNTHESIZED_WIRE_1589));


OneBitAdder	b2v_inst617(
	.ci(SYNTHESIZED_WIRE_1697),
	.a(SYNTHESIZED_WIRE_1698),
	.b(SYNTHESIZED_WIRE_1699),
	.co(SYNTHESIZED_WIRE_1700),
	.s(SYNTHESIZED_WIRE_1592));


OneBitAdder	b2v_inst618(
	.ci(SYNTHESIZED_WIRE_1700),
	.a(SYNTHESIZED_WIRE_1701),
	.b(SYNTHESIZED_WIRE_1702),
	.co(SYNTHESIZED_WIRE_1703),
	.s(SYNTHESIZED_WIRE_1595));


OneBitAdder	b2v_inst619(
	.ci(SYNTHESIZED_WIRE_1703),
	.a(SYNTHESIZED_WIRE_1704),
	.b(SYNTHESIZED_WIRE_1705),
	.co(SYNTHESIZED_WIRE_1709),
	.s(SYNTHESIZED_WIRE_1598));


OneBitAdder	b2v_inst62(
	.ci(SYNTHESIZED_WIRE_1706),
	.a(SYNTHESIZED_WIRE_1707),
	.b(SYNTHESIZED_WIRE_1708),
	.co(SYNTHESIZED_WIRE_1739),
	.s(Z_ALTERA_SYNTHESIZED[44]));


OneBitAdder	b2v_inst620(
	.ci(SYNTHESIZED_WIRE_1709),
	.a(SYNTHESIZED_WIRE_1710),
	.b(SYNTHESIZED_WIRE_1711),
	.co(SYNTHESIZED_WIRE_1712),
	.s(SYNTHESIZED_WIRE_1601));


OneBitAdder	b2v_inst621(
	.ci(SYNTHESIZED_WIRE_1712),
	.a(SYNTHESIZED_WIRE_1713),
	.b(SYNTHESIZED_WIRE_1714),
	.co(SYNTHESIZED_WIRE_1715),
	.s(SYNTHESIZED_WIRE_1604));


OneBitAdder	b2v_inst622(
	.ci(SYNTHESIZED_WIRE_1715),
	.a(SYNTHESIZED_WIRE_1716),
	.b(SYNTHESIZED_WIRE_1717),
	.co(SYNTHESIZED_WIRE_1718),
	.s(SYNTHESIZED_WIRE_1607));


OneBitAdder	b2v_inst623(
	.ci(SYNTHESIZED_WIRE_1718),
	.a(SYNTHESIZED_WIRE_1719),
	.b(SYNTHESIZED_WIRE_1720),
	.co(SYNTHESIZED_WIRE_1721),
	.s(SYNTHESIZED_WIRE_1613));


OneBitAdder	b2v_inst624(
	.ci(SYNTHESIZED_WIRE_1721),
	.a(SYNTHESIZED_WIRE_1722),
	.b(SYNTHESIZED_WIRE_1723),
	.co(SYNTHESIZED_WIRE_1619),
	.s(SYNTHESIZED_WIRE_1616));


OneBitAdder	b2v_inst625(
	.ci(SYNTHESIZED_WIRE_1724),
	.a(SYNTHESIZED_WIRE_1725),
	.b(SYNTHESIZED_WIRE_1726),
	.co(SYNTHESIZED_WIRE_1727),
	.s(SYNTHESIZED_WIRE_1567));


OneBitAdder	b2v_inst626(
	.ci(SYNTHESIZED_WIRE_1727),
	.a(SYNTHESIZED_WIRE_1728),
	.b(SYNTHESIZED_WIRE_1729),
	.co(SYNTHESIZED_WIRE_1730),
	.s(SYNTHESIZED_WIRE_1622));


OneBitAdder	b2v_inst627(
	.ci(SYNTHESIZED_WIRE_1730),
	.a(SYNTHESIZED_WIRE_1731),
	.b(SYNTHESIZED_WIRE_1732),
	.co(SYNTHESIZED_WIRE_1733),
	.s(SYNTHESIZED_WIRE_1625));


OneBitAdder	b2v_inst628(
	.ci(SYNTHESIZED_WIRE_1733),
	.a(SYNTHESIZED_WIRE_1734),
	.b(SYNTHESIZED_WIRE_1735),
	.co(SYNTHESIZED_WIRE_1736),
	.s(SYNTHESIZED_WIRE_1628));


OneBitAdder	b2v_inst629(
	.ci(SYNTHESIZED_WIRE_1736),
	.a(SYNTHESIZED_WIRE_1737),
	.b(SYNTHESIZED_WIRE_1738),
	.co(SYNTHESIZED_WIRE_1742),
	.s(SYNTHESIZED_WIRE_1631));


OneBitAdder	b2v_inst63(
	.ci(SYNTHESIZED_WIRE_1739),
	.a(SYNTHESIZED_WIRE_1740),
	.b(SYNTHESIZED_WIRE_1741),
	.co(SYNTHESIZED_WIRE_1772),
	.s(Z_ALTERA_SYNTHESIZED[45]));


OneBitAdder	b2v_inst630(
	.ci(SYNTHESIZED_WIRE_1742),
	.a(SYNTHESIZED_WIRE_1743),
	.b(SYNTHESIZED_WIRE_1744),
	.co(SYNTHESIZED_WIRE_1745),
	.s(SYNTHESIZED_WIRE_1634));


OneBitAdder	b2v_inst631(
	.ci(SYNTHESIZED_WIRE_1745),
	.a(SYNTHESIZED_WIRE_1746),
	.b(SYNTHESIZED_WIRE_1747),
	.co(SYNTHESIZED_WIRE_1748),
	.s(SYNTHESIZED_WIRE_1637));


OneBitAdder	b2v_inst632(
	.ci(SYNTHESIZED_WIRE_1748),
	.a(SYNTHESIZED_WIRE_1749),
	.b(SYNTHESIZED_WIRE_1750),
	.co(SYNTHESIZED_WIRE_1751),
	.s(SYNTHESIZED_WIRE_1640));


OneBitAdder	b2v_inst633(
	.ci(SYNTHESIZED_WIRE_1751),
	.a(SYNTHESIZED_WIRE_1752),
	.b(SYNTHESIZED_WIRE_1753),
	.co(SYNTHESIZED_WIRE_1754),
	.s(SYNTHESIZED_WIRE_1646));


OneBitAdder	b2v_inst634(
	.ci(SYNTHESIZED_WIRE_1754),
	.a(SYNTHESIZED_WIRE_1755),
	.b(SYNTHESIZED_WIRE_1756),
	.co(SYNTHESIZED_WIRE_1757),
	.s(SYNTHESIZED_WIRE_1649));


OneBitAdder	b2v_inst635(
	.ci(SYNTHESIZED_WIRE_1757),
	.a(SYNTHESIZED_WIRE_1758),
	.b(SYNTHESIZED_WIRE_1759),
	.co(SYNTHESIZED_WIRE_1760),
	.s(SYNTHESIZED_WIRE_1652));


OneBitAdder	b2v_inst636(
	.ci(SYNTHESIZED_WIRE_1760),
	.a(SYNTHESIZED_WIRE_1761),
	.b(SYNTHESIZED_WIRE_1762),
	.co(SYNTHESIZED_WIRE_1763),
	.s(SYNTHESIZED_WIRE_1655));


OneBitAdder	b2v_inst637(
	.ci(SYNTHESIZED_WIRE_1763),
	.a(SYNTHESIZED_WIRE_1764),
	.b(SYNTHESIZED_WIRE_1765),
	.co(SYNTHESIZED_WIRE_1766),
	.s(SYNTHESIZED_WIRE_1658));


OneBitAdder	b2v_inst638(
	.ci(SYNTHESIZED_WIRE_1766),
	.a(SYNTHESIZED_WIRE_1767),
	.b(SYNTHESIZED_WIRE_1768),
	.co(SYNTHESIZED_WIRE_1769),
	.s(SYNTHESIZED_WIRE_1661));


OneBitAdder	b2v_inst639(
	.ci(SYNTHESIZED_WIRE_1769),
	.a(SYNTHESIZED_WIRE_1770),
	.b(SYNTHESIZED_WIRE_1771),
	.co(SYNTHESIZED_WIRE_1775),
	.s(SYNTHESIZED_WIRE_1664));


OneBitAdder	b2v_inst64(
	.ci(SYNTHESIZED_WIRE_1772),
	.a(SYNTHESIZED_WIRE_1773),
	.b(SYNTHESIZED_WIRE_1774),
	.co(SYNTHESIZED_WIRE_1804),
	.s(Z_ALTERA_SYNTHESIZED[46]));


OneBitAdder	b2v_inst640(
	.ci(SYNTHESIZED_WIRE_1775),
	.a(SYNTHESIZED_WIRE_1776),
	.b(SYNTHESIZED_WIRE_1777),
	.co(SYNTHESIZED_WIRE_1676),
	.s(SYNTHESIZED_WIRE_1667));


OneBitAdderHalf	b2v_inst641(
	.A(SYNTHESIZED_WIRE_1778),
	.B(SYNTHESIZED_WIRE_1779),
	.C(SYNTHESIZED_WIRE_1828),
	.S(Z_ALTERA_SYNTHESIZED[12]));


OneBitAdder	b2v_inst642(
	.ci(SYNTHESIZED_WIRE_1780),
	.a(SYNTHESIZED_WIRE_1781),
	.b(SYNTHESIZED_WIRE_1782),
	.co(SYNTHESIZED_WIRE_1783),
	.s(SYNTHESIZED_WIRE_1777));


OneBitAdder	b2v_inst643(
	.ci(SYNTHESIZED_WIRE_1783),
	.a(SYNTHESIZED_WIRE_1784),
	.b(SYNTHESIZED_WIRE_1785),
	.co(SYNTHESIZED_WIRE_1786),
	.s(SYNTHESIZED_WIRE_1678));


OneBitAdder	b2v_inst644(
	.ci(SYNTHESIZED_WIRE_1786),
	.a(SYNTHESIZED_WIRE_1787),
	.b(SYNTHESIZED_WIRE_1788),
	.co(SYNTHESIZED_WIRE_1789),
	.s(SYNTHESIZED_WIRE_1681));


OneBitAdder	b2v_inst645(
	.ci(SYNTHESIZED_WIRE_1789),
	.a(SYNTHESIZED_WIRE_1790),
	.b(SYNTHESIZED_WIRE_1791),
	.co(SYNTHESIZED_WIRE_1792),
	.s(SYNTHESIZED_WIRE_1684));


OneBitAdder	b2v_inst646(
	.ci(SYNTHESIZED_WIRE_1792),
	.a(SYNTHESIZED_WIRE_1793),
	.b(SYNTHESIZED_WIRE_1794),
	.co(SYNTHESIZED_WIRE_1795),
	.s(SYNTHESIZED_WIRE_1687));


OneBitAdder	b2v_inst647(
	.ci(SYNTHESIZED_WIRE_1795),
	.a(SYNTHESIZED_WIRE_1796),
	.b(SYNTHESIZED_WIRE_1797),
	.co(SYNTHESIZED_WIRE_1798),
	.s(SYNTHESIZED_WIRE_1690));


OneBitAdder	b2v_inst648(
	.ci(SYNTHESIZED_WIRE_1798),
	.a(SYNTHESIZED_WIRE_1799),
	.b(SYNTHESIZED_WIRE_1800),
	.co(SYNTHESIZED_WIRE_1801),
	.s(SYNTHESIZED_WIRE_1693));


OneBitAdder	b2v_inst649(
	.ci(SYNTHESIZED_WIRE_1801),
	.a(SYNTHESIZED_WIRE_1802),
	.b(SYNTHESIZED_WIRE_1803),
	.co(SYNTHESIZED_WIRE_1807),
	.s(SYNTHESIZED_WIRE_1696));


OneBitAdder	b2v_inst65(
	.ci(SYNTHESIZED_WIRE_1804),
	.a(SYNTHESIZED_WIRE_1805),
	.b(SYNTHESIZED_WIRE_1806),
	.co(SYNTHESIZED_WIRE_824),
	.s(Z_ALTERA_SYNTHESIZED[47]));


OneBitAdder	b2v_inst650(
	.ci(SYNTHESIZED_WIRE_1807),
	.a(SYNTHESIZED_WIRE_1808),
	.b(SYNTHESIZED_WIRE_1809),
	.co(SYNTHESIZED_WIRE_1810),
	.s(SYNTHESIZED_WIRE_1699));


OneBitAdder	b2v_inst651(
	.ci(SYNTHESIZED_WIRE_1810),
	.a(SYNTHESIZED_WIRE_1811),
	.b(SYNTHESIZED_WIRE_1812),
	.co(SYNTHESIZED_WIRE_1813),
	.s(SYNTHESIZED_WIRE_1702));


OneBitAdder	b2v_inst652(
	.ci(SYNTHESIZED_WIRE_1813),
	.a(SYNTHESIZED_WIRE_1814),
	.b(SYNTHESIZED_WIRE_1815),
	.co(SYNTHESIZED_WIRE_1816),
	.s(SYNTHESIZED_WIRE_1705));


OneBitAdder	b2v_inst653(
	.ci(SYNTHESIZED_WIRE_1816),
	.a(SYNTHESIZED_WIRE_1817),
	.b(SYNTHESIZED_WIRE_1818),
	.co(SYNTHESIZED_WIRE_1819),
	.s(SYNTHESIZED_WIRE_1711));


OneBitAdder	b2v_inst654(
	.ci(SYNTHESIZED_WIRE_1819),
	.a(SYNTHESIZED_WIRE_1820),
	.b(SYNTHESIZED_WIRE_1821),
	.co(SYNTHESIZED_WIRE_1822),
	.s(SYNTHESIZED_WIRE_1714));


OneBitAdder	b2v_inst655(
	.ci(SYNTHESIZED_WIRE_1822),
	.a(SYNTHESIZED_WIRE_1823),
	.b(SYNTHESIZED_WIRE_1824),
	.co(SYNTHESIZED_WIRE_1825),
	.s(SYNTHESIZED_WIRE_1717));


OneBitAdder	b2v_inst656(
	.ci(SYNTHESIZED_WIRE_1825),
	.a(SYNTHESIZED_WIRE_1826),
	.b(SYNTHESIZED_WIRE_1827),
	.co(SYNTHESIZED_WIRE_1723),
	.s(SYNTHESIZED_WIRE_1720));


OneBitAdder	b2v_inst657(
	.ci(SYNTHESIZED_WIRE_1828),
	.a(SYNTHESIZED_WIRE_1829),
	.b(SYNTHESIZED_WIRE_1830),
	.co(SYNTHESIZED_WIRE_1831),
	.s(SYNTHESIZED_WIRE_1671));


OneBitAdder	b2v_inst658(
	.ci(SYNTHESIZED_WIRE_1831),
	.a(SYNTHESIZED_WIRE_1832),
	.b(SYNTHESIZED_WIRE_1833),
	.co(SYNTHESIZED_WIRE_1834),
	.s(SYNTHESIZED_WIRE_1726));


OneBitAdder	b2v_inst659(
	.ci(SYNTHESIZED_WIRE_1834),
	.a(SYNTHESIZED_WIRE_1835),
	.b(SYNTHESIZED_WIRE_1836),
	.co(SYNTHESIZED_WIRE_1840),
	.s(SYNTHESIZED_WIRE_1729));


OneBitAdder	b2v_inst66(
	.ci(SYNTHESIZED_WIRE_1837),
	.a(SYNTHESIZED_WIRE_1838),
	.b(SYNTHESIZED_WIRE_1839),
	.co(SYNTHESIZED_WIRE_1870),
	.s(SYNTHESIZED_WIRE_1806));


OneBitAdder	b2v_inst660(
	.ci(SYNTHESIZED_WIRE_1840),
	.a(SYNTHESIZED_WIRE_1841),
	.b(SYNTHESIZED_WIRE_1842),
	.co(SYNTHESIZED_WIRE_1843),
	.s(SYNTHESIZED_WIRE_1732));


OneBitAdder	b2v_inst661(
	.ci(SYNTHESIZED_WIRE_1843),
	.a(SYNTHESIZED_WIRE_1844),
	.b(SYNTHESIZED_WIRE_1845),
	.co(SYNTHESIZED_WIRE_1846),
	.s(SYNTHESIZED_WIRE_1735));


OneBitAdder	b2v_inst662(
	.ci(SYNTHESIZED_WIRE_1846),
	.a(SYNTHESIZED_WIRE_1847),
	.b(SYNTHESIZED_WIRE_1848),
	.co(SYNTHESIZED_WIRE_1849),
	.s(SYNTHESIZED_WIRE_1738));


OneBitAdder	b2v_inst663(
	.ci(SYNTHESIZED_WIRE_1849),
	.a(SYNTHESIZED_WIRE_1850),
	.b(SYNTHESIZED_WIRE_1851),
	.co(SYNTHESIZED_WIRE_1852),
	.s(SYNTHESIZED_WIRE_1744));


OneBitAdder	b2v_inst664(
	.ci(SYNTHESIZED_WIRE_1852),
	.a(SYNTHESIZED_WIRE_1853),
	.b(SYNTHESIZED_WIRE_1854),
	.co(SYNTHESIZED_WIRE_1855),
	.s(SYNTHESIZED_WIRE_1747));


OneBitAdder	b2v_inst665(
	.ci(SYNTHESIZED_WIRE_1855),
	.a(SYNTHESIZED_WIRE_1856),
	.b(SYNTHESIZED_WIRE_1857),
	.co(SYNTHESIZED_WIRE_1858),
	.s(SYNTHESIZED_WIRE_1750));


OneBitAdder	b2v_inst666(
	.ci(SYNTHESIZED_WIRE_1858),
	.a(SYNTHESIZED_WIRE_1859),
	.b(SYNTHESIZED_WIRE_1860),
	.co(SYNTHESIZED_WIRE_1861),
	.s(SYNTHESIZED_WIRE_1753));


OneBitAdder	b2v_inst667(
	.ci(SYNTHESIZED_WIRE_1861),
	.a(SYNTHESIZED_WIRE_1862),
	.b(SYNTHESIZED_WIRE_1863),
	.co(SYNTHESIZED_WIRE_1864),
	.s(SYNTHESIZED_WIRE_1756));


OneBitAdder	b2v_inst668(
	.ci(SYNTHESIZED_WIRE_1864),
	.a(SYNTHESIZED_WIRE_1865),
	.b(SYNTHESIZED_WIRE_1866),
	.co(SYNTHESIZED_WIRE_1867),
	.s(SYNTHESIZED_WIRE_1759));


OneBitAdder	b2v_inst669(
	.ci(SYNTHESIZED_WIRE_1867),
	.a(SYNTHESIZED_WIRE_1868),
	.b(SYNTHESIZED_WIRE_1869),
	.co(SYNTHESIZED_WIRE_1873),
	.s(SYNTHESIZED_WIRE_1762));


OneBitAdder	b2v_inst67(
	.ci(SYNTHESIZED_WIRE_1870),
	.a(SYNTHESIZED_WIRE_1871),
	.b(SYNTHESIZED_WIRE_1872),
	.co(SYNTHESIZED_WIRE_1902),
	.s(SYNTHESIZED_WIRE_826));


OneBitAdder	b2v_inst670(
	.ci(SYNTHESIZED_WIRE_1873),
	.a(SYNTHESIZED_WIRE_1874),
	.b(SYNTHESIZED_WIRE_1875),
	.co(SYNTHESIZED_WIRE_1876),
	.s(SYNTHESIZED_WIRE_1765));


OneBitAdder	b2v_inst671(
	.ci(SYNTHESIZED_WIRE_1876),
	.a(SYNTHESIZED_WIRE_1877),
	.b(SYNTHESIZED_WIRE_1878),
	.co(SYNTHESIZED_WIRE_1879),
	.s(SYNTHESIZED_WIRE_1768));


OneBitAdder	b2v_inst672(
	.ci(SYNTHESIZED_WIRE_1879),
	.a(SYNTHESIZED_WIRE_1880),
	.b(SYNTHESIZED_WIRE_1881),
	.co(SYNTHESIZED_WIRE_1780),
	.s(SYNTHESIZED_WIRE_1771));


OneBitAdderHalf	b2v_inst673(
	.A(SYNTHESIZED_WIRE_1882),
	.B(SYNTHESIZED_WIRE_1883),
	.C(SYNTHESIZED_WIRE_1932),
	.S(Z_ALTERA_SYNTHESIZED[11]));


OneBitAdder	b2v_inst674(
	.ci(SYNTHESIZED_WIRE_1884),
	.a(SYNTHESIZED_WIRE_1885),
	.b(SYNTHESIZED_WIRE_1886),
	.co(SYNTHESIZED_WIRE_1887),
	.s(SYNTHESIZED_WIRE_1881));


OneBitAdder	b2v_inst675(
	.ci(SYNTHESIZED_WIRE_1887),
	.a(SYNTHESIZED_WIRE_1888),
	.b(SYNTHESIZED_WIRE_1889),
	.co(SYNTHESIZED_WIRE_1890),
	.s(SYNTHESIZED_WIRE_1782));


OneBitAdder	b2v_inst676(
	.ci(SYNTHESIZED_WIRE_1890),
	.a(SYNTHESIZED_WIRE_1891),
	.b(SYNTHESIZED_WIRE_1892),
	.co(SYNTHESIZED_WIRE_1893),
	.s(SYNTHESIZED_WIRE_1785));


OneBitAdder	b2v_inst677(
	.ci(SYNTHESIZED_WIRE_1893),
	.a(SYNTHESIZED_WIRE_1894),
	.b(SYNTHESIZED_WIRE_1895),
	.co(SYNTHESIZED_WIRE_1896),
	.s(SYNTHESIZED_WIRE_1788));


OneBitAdder	b2v_inst678(
	.ci(SYNTHESIZED_WIRE_1896),
	.a(SYNTHESIZED_WIRE_1897),
	.b(SYNTHESIZED_WIRE_1898),
	.co(SYNTHESIZED_WIRE_1899),
	.s(SYNTHESIZED_WIRE_1791));


OneBitAdder	b2v_inst679(
	.ci(SYNTHESIZED_WIRE_1899),
	.a(SYNTHESIZED_WIRE_1900),
	.b(SYNTHESIZED_WIRE_1901),
	.co(SYNTHESIZED_WIRE_1905),
	.s(SYNTHESIZED_WIRE_1794));


OneBitAdder	b2v_inst68(
	.ci(SYNTHESIZED_WIRE_1902),
	.a(SYNTHESIZED_WIRE_1903),
	.b(SYNTHESIZED_WIRE_1904),
	.co(SYNTHESIZED_WIRE_1935),
	.s(SYNTHESIZED_WIRE_858));


OneBitAdder	b2v_inst680(
	.ci(SYNTHESIZED_WIRE_1905),
	.a(SYNTHESIZED_WIRE_1906),
	.b(SYNTHESIZED_WIRE_1907),
	.co(SYNTHESIZED_WIRE_1908),
	.s(SYNTHESIZED_WIRE_1797));


OneBitAdder	b2v_inst681(
	.ci(SYNTHESIZED_WIRE_1908),
	.a(SYNTHESIZED_WIRE_1909),
	.b(SYNTHESIZED_WIRE_1910),
	.co(SYNTHESIZED_WIRE_1911),
	.s(SYNTHESIZED_WIRE_1800));


OneBitAdder	b2v_inst682(
	.ci(SYNTHESIZED_WIRE_1911),
	.a(SYNTHESIZED_WIRE_1912),
	.b(SYNTHESIZED_WIRE_1913),
	.co(SYNTHESIZED_WIRE_1914),
	.s(SYNTHESIZED_WIRE_1803));


OneBitAdder	b2v_inst683(
	.ci(SYNTHESIZED_WIRE_1914),
	.a(SYNTHESIZED_WIRE_1915),
	.b(SYNTHESIZED_WIRE_1916),
	.co(SYNTHESIZED_WIRE_1917),
	.s(SYNTHESIZED_WIRE_1809));


OneBitAdder	b2v_inst684(
	.ci(SYNTHESIZED_WIRE_1917),
	.a(SYNTHESIZED_WIRE_1918),
	.b(SYNTHESIZED_WIRE_1919),
	.co(SYNTHESIZED_WIRE_1920),
	.s(SYNTHESIZED_WIRE_1812));


OneBitAdder	b2v_inst685(
	.ci(SYNTHESIZED_WIRE_1920),
	.a(SYNTHESIZED_WIRE_1921),
	.b(SYNTHESIZED_WIRE_1922),
	.co(SYNTHESIZED_WIRE_1923),
	.s(SYNTHESIZED_WIRE_1815));


OneBitAdder	b2v_inst686(
	.ci(SYNTHESIZED_WIRE_1923),
	.a(SYNTHESIZED_WIRE_1924),
	.b(SYNTHESIZED_WIRE_1925),
	.co(SYNTHESIZED_WIRE_1926),
	.s(SYNTHESIZED_WIRE_1818));


OneBitAdder	b2v_inst687(
	.ci(SYNTHESIZED_WIRE_1926),
	.a(SYNTHESIZED_WIRE_1927),
	.b(SYNTHESIZED_WIRE_1928),
	.co(SYNTHESIZED_WIRE_1929),
	.s(SYNTHESIZED_WIRE_1821));


OneBitAdder	b2v_inst688(
	.ci(SYNTHESIZED_WIRE_1929),
	.a(SYNTHESIZED_WIRE_1930),
	.b(SYNTHESIZED_WIRE_1931),
	.co(SYNTHESIZED_WIRE_1827),
	.s(SYNTHESIZED_WIRE_1824));


OneBitAdder	b2v_inst689(
	.ci(SYNTHESIZED_WIRE_1932),
	.a(SYNTHESIZED_WIRE_1933),
	.b(SYNTHESIZED_WIRE_1934),
	.co(SYNTHESIZED_WIRE_1938),
	.s(SYNTHESIZED_WIRE_1778));


OneBitAdder	b2v_inst69(
	.ci(SYNTHESIZED_WIRE_1935),
	.a(SYNTHESIZED_WIRE_1936),
	.b(SYNTHESIZED_WIRE_1937),
	.co(SYNTHESIZED_WIRE_1968),
	.s(SYNTHESIZED_WIRE_891));


OneBitAdder	b2v_inst690(
	.ci(SYNTHESIZED_WIRE_1938),
	.a(SYNTHESIZED_WIRE_1939),
	.b(SYNTHESIZED_WIRE_1940),
	.co(SYNTHESIZED_WIRE_1941),
	.s(SYNTHESIZED_WIRE_1830));


OneBitAdder	b2v_inst691(
	.ci(SYNTHESIZED_WIRE_1941),
	.a(SYNTHESIZED_WIRE_1942),
	.b(SYNTHESIZED_WIRE_1943),
	.co(SYNTHESIZED_WIRE_1944),
	.s(SYNTHESIZED_WIRE_1833));


OneBitAdder	b2v_inst692(
	.ci(SYNTHESIZED_WIRE_1944),
	.a(SYNTHESIZED_WIRE_1945),
	.b(SYNTHESIZED_WIRE_1946),
	.co(SYNTHESIZED_WIRE_1947),
	.s(SYNTHESIZED_WIRE_1836));


OneBitAdder	b2v_inst693(
	.ci(SYNTHESIZED_WIRE_1947),
	.a(SYNTHESIZED_WIRE_1948),
	.b(SYNTHESIZED_WIRE_1949),
	.co(SYNTHESIZED_WIRE_1950),
	.s(SYNTHESIZED_WIRE_1842));


OneBitAdder	b2v_inst694(
	.ci(SYNTHESIZED_WIRE_1950),
	.a(SYNTHESIZED_WIRE_1951),
	.b(SYNTHESIZED_WIRE_1952),
	.co(SYNTHESIZED_WIRE_1953),
	.s(SYNTHESIZED_WIRE_1845));


OneBitAdder	b2v_inst695(
	.ci(SYNTHESIZED_WIRE_1953),
	.a(SYNTHESIZED_WIRE_1954),
	.b(SYNTHESIZED_WIRE_1955),
	.co(SYNTHESIZED_WIRE_1956),
	.s(SYNTHESIZED_WIRE_1848));


OneBitAdder	b2v_inst696(
	.ci(SYNTHESIZED_WIRE_1956),
	.a(SYNTHESIZED_WIRE_1957),
	.b(SYNTHESIZED_WIRE_1958),
	.co(SYNTHESIZED_WIRE_1959),
	.s(SYNTHESIZED_WIRE_1851));


OneBitAdder	b2v_inst697(
	.ci(SYNTHESIZED_WIRE_1959),
	.a(SYNTHESIZED_WIRE_1960),
	.b(SYNTHESIZED_WIRE_1961),
	.co(SYNTHESIZED_WIRE_1962),
	.s(SYNTHESIZED_WIRE_1854));


OneBitAdder	b2v_inst698(
	.ci(SYNTHESIZED_WIRE_1962),
	.a(SYNTHESIZED_WIRE_1963),
	.b(SYNTHESIZED_WIRE_1964),
	.co(SYNTHESIZED_WIRE_1965),
	.s(SYNTHESIZED_WIRE_1857));


OneBitAdder	b2v_inst699(
	.ci(SYNTHESIZED_WIRE_1965),
	.a(SYNTHESIZED_WIRE_1966),
	.b(SYNTHESIZED_WIRE_1967),
	.co(SYNTHESIZED_WIRE_1971),
	.s(SYNTHESIZED_WIRE_1860));


OneBitAdder	b2v_inst70(
	.ci(SYNTHESIZED_WIRE_1968),
	.a(SYNTHESIZED_WIRE_1969),
	.b(SYNTHESIZED_WIRE_1970),
	.co(SYNTHESIZED_WIRE_2000),
	.s(SYNTHESIZED_WIRE_924));


OneBitAdder	b2v_inst700(
	.ci(SYNTHESIZED_WIRE_1971),
	.a(SYNTHESIZED_WIRE_1972),
	.b(SYNTHESIZED_WIRE_1973),
	.co(SYNTHESIZED_WIRE_1974),
	.s(SYNTHESIZED_WIRE_1863));


OneBitAdder	b2v_inst701(
	.ci(SYNTHESIZED_WIRE_1974),
	.a(SYNTHESIZED_WIRE_1975),
	.b(SYNTHESIZED_WIRE_1976),
	.co(SYNTHESIZED_WIRE_1977),
	.s(SYNTHESIZED_WIRE_1866));


OneBitAdder	b2v_inst702(
	.ci(SYNTHESIZED_WIRE_1977),
	.a(SYNTHESIZED_WIRE_1978),
	.b(SYNTHESIZED_WIRE_1979),
	.co(SYNTHESIZED_WIRE_1980),
	.s(SYNTHESIZED_WIRE_1869));


OneBitAdder	b2v_inst703(
	.ci(SYNTHESIZED_WIRE_1980),
	.a(SYNTHESIZED_WIRE_1981),
	.b(SYNTHESIZED_WIRE_1982),
	.co(SYNTHESIZED_WIRE_1983),
	.s(SYNTHESIZED_WIRE_1875));


OneBitAdder	b2v_inst704(
	.ci(SYNTHESIZED_WIRE_1983),
	.a(SYNTHESIZED_WIRE_1984),
	.b(SYNTHESIZED_WIRE_1985),
	.co(SYNTHESIZED_WIRE_1884),
	.s(SYNTHESIZED_WIRE_1878));


OneBitAdderHalf	b2v_inst705(
	.A(SYNTHESIZED_WIRE_1986),
	.B(SYNTHESIZED_WIRE_1987),
	.C(SYNTHESIZED_WIRE_2039),
	.S(Z_ALTERA_SYNTHESIZED[10]));


OneBitAdder	b2v_inst706(
	.ci(SYNTHESIZED_WIRE_1988),
	.a(SYNTHESIZED_WIRE_1989),
	.b(SYNTHESIZED_WIRE_1990),
	.co(SYNTHESIZED_WIRE_1991),
	.s(SYNTHESIZED_WIRE_1985));


OneBitAdder	b2v_inst707(
	.ci(SYNTHESIZED_WIRE_1991),
	.a(SYNTHESIZED_WIRE_1992),
	.b(SYNTHESIZED_WIRE_1993),
	.co(SYNTHESIZED_WIRE_1994),
	.s(SYNTHESIZED_WIRE_1886));


OneBitAdder	b2v_inst708(
	.ci(SYNTHESIZED_WIRE_1994),
	.a(SYNTHESIZED_WIRE_1995),
	.b(SYNTHESIZED_WIRE_1996),
	.co(SYNTHESIZED_WIRE_1997),
	.s(SYNTHESIZED_WIRE_1889));


OneBitAdder	b2v_inst709(
	.ci(SYNTHESIZED_WIRE_1997),
	.a(SYNTHESIZED_WIRE_1998),
	.b(SYNTHESIZED_WIRE_1999),
	.co(SYNTHESIZED_WIRE_2003),
	.s(SYNTHESIZED_WIRE_1892));


OneBitAdder	b2v_inst71(
	.ci(SYNTHESIZED_WIRE_2000),
	.a(SYNTHESIZED_WIRE_2001),
	.b(SYNTHESIZED_WIRE_2002),
	.co(SYNTHESIZED_WIRE_2033),
	.s(SYNTHESIZED_WIRE_956));


OneBitAdder	b2v_inst710(
	.ci(SYNTHESIZED_WIRE_2003),
	.a(SYNTHESIZED_WIRE_2004),
	.b(SYNTHESIZED_WIRE_2005),
	.co(SYNTHESIZED_WIRE_2006),
	.s(SYNTHESIZED_WIRE_1895));


OneBitAdder	b2v_inst711(
	.ci(SYNTHESIZED_WIRE_2006),
	.a(SYNTHESIZED_WIRE_2007),
	.b(SYNTHESIZED_WIRE_2008),
	.co(SYNTHESIZED_WIRE_2009),
	.s(SYNTHESIZED_WIRE_1898));


OneBitAdder	b2v_inst712(
	.ci(SYNTHESIZED_WIRE_2009),
	.a(SYNTHESIZED_WIRE_2010),
	.b(SYNTHESIZED_WIRE_2011),
	.co(SYNTHESIZED_WIRE_2012),
	.s(SYNTHESIZED_WIRE_1901));


OneBitAdder	b2v_inst713(
	.ci(SYNTHESIZED_WIRE_2012),
	.a(SYNTHESIZED_WIRE_2013),
	.b(SYNTHESIZED_WIRE_2014),
	.co(SYNTHESIZED_WIRE_2015),
	.s(SYNTHESIZED_WIRE_1907));


OneBitAdder	b2v_inst714(
	.ci(SYNTHESIZED_WIRE_2015),
	.a(SYNTHESIZED_WIRE_2016),
	.b(SYNTHESIZED_WIRE_2017),
	.co(SYNTHESIZED_WIRE_2018),
	.s(SYNTHESIZED_WIRE_1910));


OneBitAdder	b2v_inst715(
	.ci(SYNTHESIZED_WIRE_2018),
	.a(SYNTHESIZED_WIRE_2019),
	.b(SYNTHESIZED_WIRE_2020),
	.co(SYNTHESIZED_WIRE_2021),
	.s(SYNTHESIZED_WIRE_1913));


OneBitAdder	b2v_inst716(
	.ci(SYNTHESIZED_WIRE_2021),
	.a(SYNTHESIZED_WIRE_2022),
	.b(SYNTHESIZED_WIRE_2023),
	.co(SYNTHESIZED_WIRE_2024),
	.s(SYNTHESIZED_WIRE_1916));


OneBitAdder	b2v_inst717(
	.ci(SYNTHESIZED_WIRE_2024),
	.a(SYNTHESIZED_WIRE_2025),
	.b(SYNTHESIZED_WIRE_2026),
	.co(SYNTHESIZED_WIRE_2027),
	.s(SYNTHESIZED_WIRE_1919));


OneBitAdder	b2v_inst718(
	.ci(SYNTHESIZED_WIRE_2027),
	.a(SYNTHESIZED_WIRE_2028),
	.b(SYNTHESIZED_WIRE_2029),
	.co(SYNTHESIZED_WIRE_2030),
	.s(SYNTHESIZED_WIRE_1922));


OneBitAdder	b2v_inst719(
	.ci(SYNTHESIZED_WIRE_2030),
	.a(SYNTHESIZED_WIRE_2031),
	.b(SYNTHESIZED_WIRE_2032),
	.co(SYNTHESIZED_WIRE_2036),
	.s(SYNTHESIZED_WIRE_1925));


OneBitAdder	b2v_inst72(
	.ci(SYNTHESIZED_WIRE_2033),
	.a(SYNTHESIZED_WIRE_2034),
	.b(SYNTHESIZED_WIRE_2035),
	.co(SYNTHESIZED_WIRE_2066),
	.s(SYNTHESIZED_WIRE_989));


OneBitAdder	b2v_inst720(
	.ci(SYNTHESIZED_WIRE_2036),
	.a(SYNTHESIZED_WIRE_2037),
	.b(SYNTHESIZED_WIRE_2038),
	.co(SYNTHESIZED_WIRE_1931),
	.s(SYNTHESIZED_WIRE_1928));


OneBitAdder	b2v_inst721(
	.ci(SYNTHESIZED_WIRE_2039),
	.a(SYNTHESIZED_WIRE_2040),
	.b(SYNTHESIZED_WIRE_2041),
	.co(SYNTHESIZED_WIRE_2042),
	.s(SYNTHESIZED_WIRE_1882));


OneBitAdder	b2v_inst722(
	.ci(SYNTHESIZED_WIRE_2042),
	.a(SYNTHESIZED_WIRE_2043),
	.b(SYNTHESIZED_WIRE_2044),
	.co(SYNTHESIZED_WIRE_2045),
	.s(SYNTHESIZED_WIRE_1934));


OneBitAdder	b2v_inst723(
	.ci(SYNTHESIZED_WIRE_2045),
	.a(SYNTHESIZED_WIRE_2046),
	.b(SYNTHESIZED_WIRE_2047),
	.co(SYNTHESIZED_WIRE_2048),
	.s(SYNTHESIZED_WIRE_1940));


OneBitAdder	b2v_inst724(
	.ci(SYNTHESIZED_WIRE_2048),
	.a(SYNTHESIZED_WIRE_2049),
	.b(SYNTHESIZED_WIRE_2050),
	.co(SYNTHESIZED_WIRE_2051),
	.s(SYNTHESIZED_WIRE_1943));


OneBitAdder	b2v_inst725(
	.ci(SYNTHESIZED_WIRE_2051),
	.a(SYNTHESIZED_WIRE_2052),
	.b(SYNTHESIZED_WIRE_2053),
	.co(SYNTHESIZED_WIRE_2054),
	.s(SYNTHESIZED_WIRE_1946));


OneBitAdder	b2v_inst726(
	.ci(SYNTHESIZED_WIRE_2054),
	.a(SYNTHESIZED_WIRE_2055),
	.b(SYNTHESIZED_WIRE_2056),
	.co(SYNTHESIZED_WIRE_2057),
	.s(SYNTHESIZED_WIRE_1949));


OneBitAdder	b2v_inst727(
	.ci(SYNTHESIZED_WIRE_2057),
	.a(SYNTHESIZED_WIRE_2058),
	.b(SYNTHESIZED_WIRE_2059),
	.co(SYNTHESIZED_WIRE_2060),
	.s(SYNTHESIZED_WIRE_1952));


OneBitAdder	b2v_inst728(
	.ci(SYNTHESIZED_WIRE_2060),
	.a(SYNTHESIZED_WIRE_2061),
	.b(SYNTHESIZED_WIRE_2062),
	.co(SYNTHESIZED_WIRE_2063),
	.s(SYNTHESIZED_WIRE_1955));


OneBitAdder	b2v_inst729(
	.ci(SYNTHESIZED_WIRE_2063),
	.a(SYNTHESIZED_WIRE_2064),
	.b(SYNTHESIZED_WIRE_2065),
	.co(SYNTHESIZED_WIRE_2069),
	.s(SYNTHESIZED_WIRE_1958));


OneBitAdder	b2v_inst73(
	.ci(SYNTHESIZED_WIRE_2066),
	.a(SYNTHESIZED_WIRE_2067),
	.b(SYNTHESIZED_WIRE_2068),
	.co(SYNTHESIZED_WIRE_2098),
	.s(SYNTHESIZED_WIRE_1022));


OneBitAdder	b2v_inst730(
	.ci(SYNTHESIZED_WIRE_2069),
	.a(SYNTHESIZED_WIRE_2070),
	.b(SYNTHESIZED_WIRE_2071),
	.co(SYNTHESIZED_WIRE_2072),
	.s(SYNTHESIZED_WIRE_1961));


OneBitAdder	b2v_inst731(
	.ci(SYNTHESIZED_WIRE_2072),
	.a(SYNTHESIZED_WIRE_2073),
	.b(SYNTHESIZED_WIRE_2074),
	.co(SYNTHESIZED_WIRE_2075),
	.s(SYNTHESIZED_WIRE_1964));


OneBitAdder	b2v_inst732(
	.ci(SYNTHESIZED_WIRE_2075),
	.a(SYNTHESIZED_WIRE_2076),
	.b(SYNTHESIZED_WIRE_2077),
	.co(SYNTHESIZED_WIRE_2078),
	.s(SYNTHESIZED_WIRE_1967));


OneBitAdder	b2v_inst733(
	.ci(SYNTHESIZED_WIRE_2078),
	.a(SYNTHESIZED_WIRE_2079),
	.b(SYNTHESIZED_WIRE_2080),
	.co(SYNTHESIZED_WIRE_2081),
	.s(SYNTHESIZED_WIRE_1973));


OneBitAdder	b2v_inst734(
	.ci(SYNTHESIZED_WIRE_2081),
	.a(SYNTHESIZED_WIRE_2082),
	.b(SYNTHESIZED_WIRE_2083),
	.co(SYNTHESIZED_WIRE_2084),
	.s(SYNTHESIZED_WIRE_1976));


OneBitAdder	b2v_inst735(
	.ci(SYNTHESIZED_WIRE_2084),
	.a(SYNTHESIZED_WIRE_2085),
	.b(SYNTHESIZED_WIRE_2086),
	.co(SYNTHESIZED_WIRE_2087),
	.s(SYNTHESIZED_WIRE_1979));


OneBitAdder	b2v_inst736(
	.ci(SYNTHESIZED_WIRE_2087),
	.a(SYNTHESIZED_WIRE_2088),
	.b(SYNTHESIZED_WIRE_2089),
	.co(SYNTHESIZED_WIRE_1988),
	.s(SYNTHESIZED_WIRE_1982));


OneBitAdderHalf	b2v_inst737(
	.A(SYNTHESIZED_WIRE_2090),
	.B(SYNTHESIZED_WIRE_2091),
	.C(SYNTHESIZED_WIRE_2143),
	.S(Z_ALTERA_SYNTHESIZED[9]));


OneBitAdder	b2v_inst738(
	.ci(SYNTHESIZED_WIRE_2092),
	.a(SYNTHESIZED_WIRE_2093),
	.b(SYNTHESIZED_WIRE_2094),
	.co(SYNTHESIZED_WIRE_2095),
	.s(SYNTHESIZED_WIRE_2089));


OneBitAdder	b2v_inst739(
	.ci(SYNTHESIZED_WIRE_2095),
	.a(SYNTHESIZED_WIRE_2096),
	.b(SYNTHESIZED_WIRE_2097),
	.co(SYNTHESIZED_WIRE_2101),
	.s(SYNTHESIZED_WIRE_1990));


OneBitAdder	b2v_inst74(
	.ci(SYNTHESIZED_WIRE_2098),
	.a(SYNTHESIZED_WIRE_2099),
	.b(SYNTHESIZED_WIRE_2100),
	.co(SYNTHESIZED_WIRE_2131),
	.s(SYNTHESIZED_WIRE_1054));


OneBitAdder	b2v_inst740(
	.ci(SYNTHESIZED_WIRE_2101),
	.a(SYNTHESIZED_WIRE_2102),
	.b(SYNTHESIZED_WIRE_2103),
	.co(SYNTHESIZED_WIRE_2104),
	.s(SYNTHESIZED_WIRE_1993));


OneBitAdder	b2v_inst741(
	.ci(SYNTHESIZED_WIRE_2104),
	.a(SYNTHESIZED_WIRE_2105),
	.b(SYNTHESIZED_WIRE_2106),
	.co(SYNTHESIZED_WIRE_2107),
	.s(SYNTHESIZED_WIRE_1996));


OneBitAdder	b2v_inst742(
	.ci(SYNTHESIZED_WIRE_2107),
	.a(SYNTHESIZED_WIRE_2108),
	.b(SYNTHESIZED_WIRE_2109),
	.co(SYNTHESIZED_WIRE_2110),
	.s(SYNTHESIZED_WIRE_1999));


OneBitAdder	b2v_inst743(
	.ci(SYNTHESIZED_WIRE_2110),
	.a(SYNTHESIZED_WIRE_2111),
	.b(SYNTHESIZED_WIRE_2112),
	.co(SYNTHESIZED_WIRE_2113),
	.s(SYNTHESIZED_WIRE_2005));


OneBitAdder	b2v_inst744(
	.ci(SYNTHESIZED_WIRE_2113),
	.a(SYNTHESIZED_WIRE_2114),
	.b(SYNTHESIZED_WIRE_2115),
	.co(SYNTHESIZED_WIRE_2116),
	.s(SYNTHESIZED_WIRE_2008));


OneBitAdder	b2v_inst745(
	.ci(SYNTHESIZED_WIRE_2116),
	.a(SYNTHESIZED_WIRE_2117),
	.b(SYNTHESIZED_WIRE_2118),
	.co(SYNTHESIZED_WIRE_2119),
	.s(SYNTHESIZED_WIRE_2011));


OneBitAdder	b2v_inst746(
	.ci(SYNTHESIZED_WIRE_2119),
	.a(SYNTHESIZED_WIRE_2120),
	.b(SYNTHESIZED_WIRE_2121),
	.co(SYNTHESIZED_WIRE_2122),
	.s(SYNTHESIZED_WIRE_2014));


OneBitAdder	b2v_inst747(
	.ci(SYNTHESIZED_WIRE_2122),
	.a(SYNTHESIZED_WIRE_2123),
	.b(SYNTHESIZED_WIRE_2124),
	.co(SYNTHESIZED_WIRE_2125),
	.s(SYNTHESIZED_WIRE_2017));


OneBitAdder	b2v_inst748(
	.ci(SYNTHESIZED_WIRE_2125),
	.a(SYNTHESIZED_WIRE_2126),
	.b(SYNTHESIZED_WIRE_2127),
	.co(SYNTHESIZED_WIRE_2128),
	.s(SYNTHESIZED_WIRE_2020));


OneBitAdder	b2v_inst749(
	.ci(SYNTHESIZED_WIRE_2128),
	.a(SYNTHESIZED_WIRE_2129),
	.b(SYNTHESIZED_WIRE_2130),
	.co(SYNTHESIZED_WIRE_2134),
	.s(SYNTHESIZED_WIRE_2023));


OneBitAdder	b2v_inst75(
	.ci(SYNTHESIZED_WIRE_2131),
	.a(SYNTHESIZED_WIRE_2132),
	.b(SYNTHESIZED_WIRE_2133),
	.co(SYNTHESIZED_WIRE_2164),
	.s(SYNTHESIZED_WIRE_1087));


OneBitAdder	b2v_inst750(
	.ci(SYNTHESIZED_WIRE_2134),
	.a(SYNTHESIZED_WIRE_2135),
	.b(SYNTHESIZED_WIRE_2136),
	.co(SYNTHESIZED_WIRE_2137),
	.s(SYNTHESIZED_WIRE_2026));


OneBitAdder	b2v_inst751(
	.ci(SYNTHESIZED_WIRE_2137),
	.a(SYNTHESIZED_WIRE_2138),
	.b(SYNTHESIZED_WIRE_2139),
	.co(SYNTHESIZED_WIRE_2140),
	.s(SYNTHESIZED_WIRE_2029));


OneBitAdder	b2v_inst752(
	.ci(SYNTHESIZED_WIRE_2140),
	.a(SYNTHESIZED_WIRE_2141),
	.b(SYNTHESIZED_WIRE_2142),
	.co(SYNTHESIZED_WIRE_2038),
	.s(SYNTHESIZED_WIRE_2032));


OneBitAdder	b2v_inst753(
	.ci(SYNTHESIZED_WIRE_2143),
	.a(SYNTHESIZED_WIRE_2144),
	.b(SYNTHESIZED_WIRE_2145),
	.co(SYNTHESIZED_WIRE_2146),
	.s(SYNTHESIZED_WIRE_1986));


OneBitAdder	b2v_inst754(
	.ci(SYNTHESIZED_WIRE_2146),
	.a(SYNTHESIZED_WIRE_2147),
	.b(SYNTHESIZED_WIRE_2148),
	.co(SYNTHESIZED_WIRE_2149),
	.s(SYNTHESIZED_WIRE_2041));


OneBitAdder	b2v_inst755(
	.ci(SYNTHESIZED_WIRE_2149),
	.a(SYNTHESIZED_WIRE_2150),
	.b(SYNTHESIZED_WIRE_2151),
	.co(SYNTHESIZED_WIRE_2152),
	.s(SYNTHESIZED_WIRE_2044));


OneBitAdder	b2v_inst756(
	.ci(SYNTHESIZED_WIRE_2152),
	.a(SYNTHESIZED_WIRE_2153),
	.b(SYNTHESIZED_WIRE_2154),
	.co(SYNTHESIZED_WIRE_2155),
	.s(SYNTHESIZED_WIRE_2047));


OneBitAdder	b2v_inst757(
	.ci(SYNTHESIZED_WIRE_2155),
	.a(SYNTHESIZED_WIRE_2156),
	.b(SYNTHESIZED_WIRE_2157),
	.co(SYNTHESIZED_WIRE_2158),
	.s(SYNTHESIZED_WIRE_2050));


OneBitAdder	b2v_inst758(
	.ci(SYNTHESIZED_WIRE_2158),
	.a(SYNTHESIZED_WIRE_2159),
	.b(SYNTHESIZED_WIRE_2160),
	.co(SYNTHESIZED_WIRE_2161),
	.s(SYNTHESIZED_WIRE_2053));


OneBitAdder	b2v_inst759(
	.ci(SYNTHESIZED_WIRE_2161),
	.a(SYNTHESIZED_WIRE_2162),
	.b(SYNTHESIZED_WIRE_2163),
	.co(SYNTHESIZED_WIRE_2167),
	.s(SYNTHESIZED_WIRE_2056));


OneBitAdder	b2v_inst76(
	.ci(SYNTHESIZED_WIRE_2164),
	.a(SYNTHESIZED_WIRE_2165),
	.b(SYNTHESIZED_WIRE_2166),
	.co(SYNTHESIZED_WIRE_2196),
	.s(SYNTHESIZED_WIRE_1120));


OneBitAdder	b2v_inst760(
	.ci(SYNTHESIZED_WIRE_2167),
	.a(SYNTHESIZED_WIRE_2168),
	.b(SYNTHESIZED_WIRE_2169),
	.co(SYNTHESIZED_WIRE_2170),
	.s(SYNTHESIZED_WIRE_2059));


OneBitAdder	b2v_inst761(
	.ci(SYNTHESIZED_WIRE_2170),
	.a(SYNTHESIZED_WIRE_2171),
	.b(SYNTHESIZED_WIRE_2172),
	.co(SYNTHESIZED_WIRE_2173),
	.s(SYNTHESIZED_WIRE_2062));


OneBitAdder	b2v_inst762(
	.ci(SYNTHESIZED_WIRE_2173),
	.a(SYNTHESIZED_WIRE_2174),
	.b(SYNTHESIZED_WIRE_2175),
	.co(SYNTHESIZED_WIRE_2176),
	.s(SYNTHESIZED_WIRE_2065));


OneBitAdder	b2v_inst763(
	.ci(SYNTHESIZED_WIRE_2176),
	.a(SYNTHESIZED_WIRE_2177),
	.b(SYNTHESIZED_WIRE_2178),
	.co(SYNTHESIZED_WIRE_2179),
	.s(SYNTHESIZED_WIRE_2071));


OneBitAdder	b2v_inst764(
	.ci(SYNTHESIZED_WIRE_2179),
	.a(SYNTHESIZED_WIRE_2180),
	.b(SYNTHESIZED_WIRE_2181),
	.co(SYNTHESIZED_WIRE_2182),
	.s(SYNTHESIZED_WIRE_2074));


OneBitAdder	b2v_inst765(
	.ci(SYNTHESIZED_WIRE_2182),
	.a(SYNTHESIZED_WIRE_2183),
	.b(SYNTHESIZED_WIRE_2184),
	.co(SYNTHESIZED_WIRE_2185),
	.s(SYNTHESIZED_WIRE_2077));


OneBitAdder	b2v_inst766(
	.ci(SYNTHESIZED_WIRE_2185),
	.a(SYNTHESIZED_WIRE_2186),
	.b(SYNTHESIZED_WIRE_2187),
	.co(SYNTHESIZED_WIRE_2188),
	.s(SYNTHESIZED_WIRE_2080));


OneBitAdder	b2v_inst767(
	.ci(SYNTHESIZED_WIRE_2188),
	.a(SYNTHESIZED_WIRE_2189),
	.b(SYNTHESIZED_WIRE_2190),
	.co(SYNTHESIZED_WIRE_2191),
	.s(SYNTHESIZED_WIRE_2083));


OneBitAdder	b2v_inst768(
	.ci(SYNTHESIZED_WIRE_2191),
	.a(SYNTHESIZED_WIRE_2192),
	.b(SYNTHESIZED_WIRE_2193),
	.co(SYNTHESIZED_WIRE_2092),
	.s(SYNTHESIZED_WIRE_2086));


OneBitAdderHalf	b2v_inst769(
	.A(SYNTHESIZED_WIRE_2194),
	.B(SYNTHESIZED_WIRE_2195),
	.C(SYNTHESIZED_WIRE_2247),
	.S(Z_ALTERA_SYNTHESIZED[8]));


OneBitAdder	b2v_inst77(
	.ci(SYNTHESIZED_WIRE_2196),
	.a(SYNTHESIZED_WIRE_2197),
	.b(SYNTHESIZED_WIRE_2198),
	.co(SYNTHESIZED_WIRE_2229),
	.s(SYNTHESIZED_WIRE_1152));


OneBitAdder	b2v_inst770(
	.ci(SYNTHESIZED_WIRE_2199),
	.a(SYNTHESIZED_WIRE_2200),
	.b(SYNTHESIZED_WIRE_2201),
	.co(SYNTHESIZED_WIRE_2202),
	.s(SYNTHESIZED_WIRE_2193));


OneBitAdder	b2v_inst771(
	.ci(SYNTHESIZED_WIRE_2202),
	.a(SYNTHESIZED_WIRE_2203),
	.b(SYNTHESIZED_WIRE_2204),
	.co(SYNTHESIZED_WIRE_2205),
	.s(SYNTHESIZED_WIRE_2094));


OneBitAdder	b2v_inst772(
	.ci(SYNTHESIZED_WIRE_2205),
	.a(SYNTHESIZED_WIRE_2206),
	.b(SYNTHESIZED_WIRE_2207),
	.co(SYNTHESIZED_WIRE_2208),
	.s(SYNTHESIZED_WIRE_2097));


OneBitAdder	b2v_inst773(
	.ci(SYNTHESIZED_WIRE_2208),
	.a(SYNTHESIZED_WIRE_2209),
	.b(SYNTHESIZED_WIRE_2210),
	.co(SYNTHESIZED_WIRE_2211),
	.s(SYNTHESIZED_WIRE_2103));


OneBitAdder	b2v_inst774(
	.ci(SYNTHESIZED_WIRE_2211),
	.a(SYNTHESIZED_WIRE_2212),
	.b(SYNTHESIZED_WIRE_2213),
	.co(SYNTHESIZED_WIRE_2214),
	.s(SYNTHESIZED_WIRE_2106));


OneBitAdder	b2v_inst775(
	.ci(SYNTHESIZED_WIRE_2214),
	.a(SYNTHESIZED_WIRE_2215),
	.b(SYNTHESIZED_WIRE_2216),
	.co(SYNTHESIZED_WIRE_2217),
	.s(SYNTHESIZED_WIRE_2109));


OneBitAdder	b2v_inst776(
	.ci(SYNTHESIZED_WIRE_2217),
	.a(SYNTHESIZED_WIRE_2218),
	.b(SYNTHESIZED_WIRE_2219),
	.co(SYNTHESIZED_WIRE_2220),
	.s(SYNTHESIZED_WIRE_2112));


OneBitAdder	b2v_inst777(
	.ci(SYNTHESIZED_WIRE_2220),
	.a(SYNTHESIZED_WIRE_2221),
	.b(SYNTHESIZED_WIRE_2222),
	.co(SYNTHESIZED_WIRE_2223),
	.s(SYNTHESIZED_WIRE_2115));


OneBitAdder	b2v_inst778(
	.ci(SYNTHESIZED_WIRE_2223),
	.a(SYNTHESIZED_WIRE_2224),
	.b(SYNTHESIZED_WIRE_2225),
	.co(SYNTHESIZED_WIRE_2226),
	.s(SYNTHESIZED_WIRE_2118));


OneBitAdder	b2v_inst779(
	.ci(SYNTHESIZED_WIRE_2226),
	.a(SYNTHESIZED_WIRE_2227),
	.b(SYNTHESIZED_WIRE_2228),
	.co(SYNTHESIZED_WIRE_2232),
	.s(SYNTHESIZED_WIRE_2121));


OneBitAdder	b2v_inst78(
	.ci(SYNTHESIZED_WIRE_2229),
	.a(SYNTHESIZED_WIRE_2230),
	.b(SYNTHESIZED_WIRE_2231),
	.co(SYNTHESIZED_WIRE_2262),
	.s(SYNTHESIZED_WIRE_1185));


OneBitAdder	b2v_inst780(
	.ci(SYNTHESIZED_WIRE_2232),
	.a(SYNTHESIZED_WIRE_2233),
	.b(SYNTHESIZED_WIRE_2234),
	.co(SYNTHESIZED_WIRE_2235),
	.s(SYNTHESIZED_WIRE_2124));


OneBitAdder	b2v_inst781(
	.ci(SYNTHESIZED_WIRE_2235),
	.a(SYNTHESIZED_WIRE_2236),
	.b(SYNTHESIZED_WIRE_2237),
	.co(SYNTHESIZED_WIRE_2238),
	.s(SYNTHESIZED_WIRE_2127));


OneBitAdder	b2v_inst782(
	.ci(SYNTHESIZED_WIRE_2238),
	.a(SYNTHESIZED_WIRE_2239),
	.b(SYNTHESIZED_WIRE_2240),
	.co(SYNTHESIZED_WIRE_2241),
	.s(SYNTHESIZED_WIRE_2130));


OneBitAdder	b2v_inst783(
	.ci(SYNTHESIZED_WIRE_2241),
	.a(SYNTHESIZED_WIRE_2242),
	.b(SYNTHESIZED_WIRE_2243),
	.co(SYNTHESIZED_WIRE_2244),
	.s(SYNTHESIZED_WIRE_2136));


OneBitAdder	b2v_inst784(
	.ci(SYNTHESIZED_WIRE_2244),
	.a(SYNTHESIZED_WIRE_2245),
	.b(SYNTHESIZED_WIRE_2246),
	.co(SYNTHESIZED_WIRE_2142),
	.s(SYNTHESIZED_WIRE_2139));


OneBitAdder	b2v_inst785(
	.ci(SYNTHESIZED_WIRE_2247),
	.a(SYNTHESIZED_WIRE_2248),
	.b(SYNTHESIZED_WIRE_2249),
	.co(SYNTHESIZED_WIRE_2250),
	.s(SYNTHESIZED_WIRE_2090));


OneBitAdder	b2v_inst786(
	.ci(SYNTHESIZED_WIRE_2250),
	.a(SYNTHESIZED_WIRE_2251),
	.b(SYNTHESIZED_WIRE_2252),
	.co(SYNTHESIZED_WIRE_2253),
	.s(SYNTHESIZED_WIRE_2145));


OneBitAdder	b2v_inst787(
	.ci(SYNTHESIZED_WIRE_2253),
	.a(SYNTHESIZED_WIRE_2254),
	.b(SYNTHESIZED_WIRE_2255),
	.co(SYNTHESIZED_WIRE_2256),
	.s(SYNTHESIZED_WIRE_2148));


OneBitAdder	b2v_inst788(
	.ci(SYNTHESIZED_WIRE_2256),
	.a(SYNTHESIZED_WIRE_2257),
	.b(SYNTHESIZED_WIRE_2258),
	.co(SYNTHESIZED_WIRE_2259),
	.s(SYNTHESIZED_WIRE_2151));


OneBitAdder	b2v_inst789(
	.ci(SYNTHESIZED_WIRE_2259),
	.a(SYNTHESIZED_WIRE_2260),
	.b(SYNTHESIZED_WIRE_2261),
	.co(SYNTHESIZED_WIRE_2265),
	.s(SYNTHESIZED_WIRE_2154));


OneBitAdder	b2v_inst79(
	.ci(SYNTHESIZED_WIRE_2262),
	.a(SYNTHESIZED_WIRE_2263),
	.b(SYNTHESIZED_WIRE_2264),
	.co(SYNTHESIZED_WIRE_2295),
	.s(SYNTHESIZED_WIRE_1218));


OneBitAdder	b2v_inst790(
	.ci(SYNTHESIZED_WIRE_2265),
	.a(SYNTHESIZED_WIRE_2266),
	.b(SYNTHESIZED_WIRE_2267),
	.co(SYNTHESIZED_WIRE_2268),
	.s(SYNTHESIZED_WIRE_2157));


OneBitAdder	b2v_inst791(
	.ci(SYNTHESIZED_WIRE_2268),
	.a(SYNTHESIZED_WIRE_2269),
	.b(SYNTHESIZED_WIRE_2270),
	.co(SYNTHESIZED_WIRE_2271),
	.s(SYNTHESIZED_WIRE_2160));


OneBitAdder	b2v_inst792(
	.ci(SYNTHESIZED_WIRE_2271),
	.a(SYNTHESIZED_WIRE_2272),
	.b(SYNTHESIZED_WIRE_2273),
	.co(SYNTHESIZED_WIRE_2274),
	.s(SYNTHESIZED_WIRE_2163));


OneBitAdder	b2v_inst793(
	.ci(SYNTHESIZED_WIRE_2274),
	.a(SYNTHESIZED_WIRE_2275),
	.b(SYNTHESIZED_WIRE_2276),
	.co(SYNTHESIZED_WIRE_2277),
	.s(SYNTHESIZED_WIRE_2169));


OneBitAdder	b2v_inst794(
	.ci(SYNTHESIZED_WIRE_2277),
	.a(SYNTHESIZED_WIRE_2278),
	.b(SYNTHESIZED_WIRE_2279),
	.co(SYNTHESIZED_WIRE_2280),
	.s(SYNTHESIZED_WIRE_2172));


OneBitAdder	b2v_inst795(
	.ci(SYNTHESIZED_WIRE_2280),
	.a(SYNTHESIZED_WIRE_2281),
	.b(SYNTHESIZED_WIRE_2282),
	.co(SYNTHESIZED_WIRE_2283),
	.s(SYNTHESIZED_WIRE_2175));


OneBitAdder	b2v_inst796(
	.ci(SYNTHESIZED_WIRE_2283),
	.a(SYNTHESIZED_WIRE_2284),
	.b(SYNTHESIZED_WIRE_2285),
	.co(SYNTHESIZED_WIRE_2286),
	.s(SYNTHESIZED_WIRE_2178));


OneBitAdder	b2v_inst797(
	.ci(SYNTHESIZED_WIRE_2286),
	.a(SYNTHESIZED_WIRE_2287),
	.b(SYNTHESIZED_WIRE_2288),
	.co(SYNTHESIZED_WIRE_2289),
	.s(SYNTHESIZED_WIRE_2181));


OneBitAdder	b2v_inst798(
	.ci(SYNTHESIZED_WIRE_2289),
	.a(SYNTHESIZED_WIRE_2290),
	.b(SYNTHESIZED_WIRE_2291),
	.co(SYNTHESIZED_WIRE_2292),
	.s(SYNTHESIZED_WIRE_2184));


OneBitAdder	b2v_inst799(
	.ci(SYNTHESIZED_WIRE_2292),
	.a(SYNTHESIZED_WIRE_2293),
	.b(SYNTHESIZED_WIRE_2294),
	.co(SYNTHESIZED_WIRE_2298),
	.s(SYNTHESIZED_WIRE_2187));


OneBitAdder	b2v_inst80(
	.ci(SYNTHESIZED_WIRE_2295),
	.a(SYNTHESIZED_WIRE_2296),
	.b(SYNTHESIZED_WIRE_2297),
	.co(SYNTHESIZED_WIRE_1283),
	.s(SYNTHESIZED_WIRE_1251));


OneBitAdder	b2v_inst800(
	.ci(SYNTHESIZED_WIRE_2298),
	.a(SYNTHESIZED_WIRE_2299),
	.b(SYNTHESIZED_WIRE_2300),
	.co(SYNTHESIZED_WIRE_2199),
	.s(SYNTHESIZED_WIRE_2190));


OneBitAdderHalf	b2v_inst801(
	.A(SYNTHESIZED_WIRE_2301),
	.B(SYNTHESIZED_WIRE_2302),
	.C(SYNTHESIZED_WIRE_2351),
	.S(Z_ALTERA_SYNTHESIZED[7]));


OneBitAdder	b2v_inst802(
	.ci(SYNTHESIZED_WIRE_2303),
	.a(SYNTHESIZED_WIRE_2304),
	.b(SYNTHESIZED_WIRE_2305),
	.co(SYNTHESIZED_WIRE_2306),
	.s(SYNTHESIZED_WIRE_2300));


OneBitAdder	b2v_inst803(
	.ci(SYNTHESIZED_WIRE_2306),
	.a(SYNTHESIZED_WIRE_2307),
	.b(SYNTHESIZED_WIRE_2308),
	.co(SYNTHESIZED_WIRE_2309),
	.s(SYNTHESIZED_WIRE_2201));


OneBitAdder	b2v_inst804(
	.ci(SYNTHESIZED_WIRE_2309),
	.a(SYNTHESIZED_WIRE_2310),
	.b(SYNTHESIZED_WIRE_2311),
	.co(SYNTHESIZED_WIRE_2312),
	.s(SYNTHESIZED_WIRE_2204));


OneBitAdder	b2v_inst805(
	.ci(SYNTHESIZED_WIRE_2312),
	.a(SYNTHESIZED_WIRE_2313),
	.b(SYNTHESIZED_WIRE_2314),
	.co(SYNTHESIZED_WIRE_2315),
	.s(SYNTHESIZED_WIRE_2207));


OneBitAdder	b2v_inst806(
	.ci(SYNTHESIZED_WIRE_2315),
	.a(SYNTHESIZED_WIRE_2316),
	.b(SYNTHESIZED_WIRE_2317),
	.co(SYNTHESIZED_WIRE_2318),
	.s(SYNTHESIZED_WIRE_2210));


OneBitAdder	b2v_inst807(
	.ci(SYNTHESIZED_WIRE_2318),
	.a(SYNTHESIZED_WIRE_2319),
	.b(SYNTHESIZED_WIRE_2320),
	.co(SYNTHESIZED_WIRE_2321),
	.s(SYNTHESIZED_WIRE_2213));


OneBitAdder	b2v_inst808(
	.ci(SYNTHESIZED_WIRE_2321),
	.a(SYNTHESIZED_WIRE_2322),
	.b(SYNTHESIZED_WIRE_2323),
	.co(SYNTHESIZED_WIRE_2324),
	.s(SYNTHESIZED_WIRE_2216));


OneBitAdder	b2v_inst809(
	.ci(SYNTHESIZED_WIRE_2324),
	.a(SYNTHESIZED_WIRE_2325),
	.b(SYNTHESIZED_WIRE_2326),
	.co(SYNTHESIZED_WIRE_2330),
	.s(SYNTHESIZED_WIRE_2219));


OneBitAdder	b2v_inst81(
	.ci(SYNTHESIZED_WIRE_2327),
	.a(SYNTHESIZED_WIRE_2328),
	.b(SYNTHESIZED_WIRE_2329),
	.co(SYNTHESIZED_WIRE_2360),
	.s(SYNTHESIZED_WIRE_0));


OneBitAdder	b2v_inst810(
	.ci(SYNTHESIZED_WIRE_2330),
	.a(SYNTHESIZED_WIRE_2331),
	.b(SYNTHESIZED_WIRE_2332),
	.co(SYNTHESIZED_WIRE_2333),
	.s(SYNTHESIZED_WIRE_2222));


OneBitAdder	b2v_inst811(
	.ci(SYNTHESIZED_WIRE_2333),
	.a(SYNTHESIZED_WIRE_2334),
	.b(SYNTHESIZED_WIRE_2335),
	.co(SYNTHESIZED_WIRE_2336),
	.s(SYNTHESIZED_WIRE_2225));


OneBitAdder	b2v_inst812(
	.ci(SYNTHESIZED_WIRE_2336),
	.a(SYNTHESIZED_WIRE_2337),
	.b(SYNTHESIZED_WIRE_2338),
	.co(SYNTHESIZED_WIRE_2339),
	.s(SYNTHESIZED_WIRE_2228));


OneBitAdder	b2v_inst813(
	.ci(SYNTHESIZED_WIRE_2339),
	.a(SYNTHESIZED_WIRE_2340),
	.b(SYNTHESIZED_WIRE_2341),
	.co(SYNTHESIZED_WIRE_2342),
	.s(SYNTHESIZED_WIRE_2234));


OneBitAdder	b2v_inst814(
	.ci(SYNTHESIZED_WIRE_2342),
	.a(SYNTHESIZED_WIRE_2343),
	.b(SYNTHESIZED_WIRE_2344),
	.co(SYNTHESIZED_WIRE_2345),
	.s(SYNTHESIZED_WIRE_2237));


OneBitAdder	b2v_inst815(
	.ci(SYNTHESIZED_WIRE_2345),
	.a(SYNTHESIZED_WIRE_2346),
	.b(SYNTHESIZED_WIRE_2347),
	.co(SYNTHESIZED_WIRE_2348),
	.s(SYNTHESIZED_WIRE_2240));


OneBitAdder	b2v_inst816(
	.ci(SYNTHESIZED_WIRE_2348),
	.a(SYNTHESIZED_WIRE_2349),
	.b(SYNTHESIZED_WIRE_2350),
	.co(SYNTHESIZED_WIRE_2246),
	.s(SYNTHESIZED_WIRE_2243));


OneBitAdder	b2v_inst817(
	.ci(SYNTHESIZED_WIRE_2351),
	.a(SYNTHESIZED_WIRE_2352),
	.b(SYNTHESIZED_WIRE_2353),
	.co(SYNTHESIZED_WIRE_2354),
	.s(SYNTHESIZED_WIRE_2194));


OneBitAdder	b2v_inst818(
	.ci(SYNTHESIZED_WIRE_2354),
	.a(SYNTHESIZED_WIRE_2355),
	.b(SYNTHESIZED_WIRE_2356),
	.co(SYNTHESIZED_WIRE_2357),
	.s(SYNTHESIZED_WIRE_2249));


OneBitAdder	b2v_inst819(
	.ci(SYNTHESIZED_WIRE_2357),
	.a(SYNTHESIZED_WIRE_2358),
	.b(SYNTHESIZED_WIRE_2359),
	.co(SYNTHESIZED_WIRE_2363),
	.s(SYNTHESIZED_WIRE_2252));


OneBitAdder	b2v_inst82(
	.ci(SYNTHESIZED_WIRE_2360),
	.a(SYNTHESIZED_WIRE_2361),
	.b(SYNTHESIZED_WIRE_2362),
	.co(SYNTHESIZED_WIRE_2393),
	.s(SYNTHESIZED_WIRE_1316));


OneBitAdder	b2v_inst820(
	.ci(SYNTHESIZED_WIRE_2363),
	.a(SYNTHESIZED_WIRE_2364),
	.b(SYNTHESIZED_WIRE_2365),
	.co(SYNTHESIZED_WIRE_2366),
	.s(SYNTHESIZED_WIRE_2255));


OneBitAdder	b2v_inst821(
	.ci(SYNTHESIZED_WIRE_2366),
	.a(SYNTHESIZED_WIRE_2367),
	.b(SYNTHESIZED_WIRE_2368),
	.co(SYNTHESIZED_WIRE_2369),
	.s(SYNTHESIZED_WIRE_2258));


OneBitAdder	b2v_inst822(
	.ci(SYNTHESIZED_WIRE_2369),
	.a(SYNTHESIZED_WIRE_2370),
	.b(SYNTHESIZED_WIRE_2371),
	.co(SYNTHESIZED_WIRE_2372),
	.s(SYNTHESIZED_WIRE_2261));


OneBitAdder	b2v_inst823(
	.ci(SYNTHESIZED_WIRE_2372),
	.a(SYNTHESIZED_WIRE_2373),
	.b(SYNTHESIZED_WIRE_2374),
	.co(SYNTHESIZED_WIRE_2375),
	.s(SYNTHESIZED_WIRE_2267));


OneBitAdder	b2v_inst824(
	.ci(SYNTHESIZED_WIRE_2375),
	.a(SYNTHESIZED_WIRE_2376),
	.b(SYNTHESIZED_WIRE_2377),
	.co(SYNTHESIZED_WIRE_2378),
	.s(SYNTHESIZED_WIRE_2270));


OneBitAdder	b2v_inst825(
	.ci(SYNTHESIZED_WIRE_2378),
	.a(SYNTHESIZED_WIRE_2379),
	.b(SYNTHESIZED_WIRE_2380),
	.co(SYNTHESIZED_WIRE_2381),
	.s(SYNTHESIZED_WIRE_2273));


OneBitAdder	b2v_inst826(
	.ci(SYNTHESIZED_WIRE_2381),
	.a(SYNTHESIZED_WIRE_2382),
	.b(SYNTHESIZED_WIRE_2383),
	.co(SYNTHESIZED_WIRE_2384),
	.s(SYNTHESIZED_WIRE_2276));


OneBitAdder	b2v_inst827(
	.ci(SYNTHESIZED_WIRE_2384),
	.a(SYNTHESIZED_WIRE_2385),
	.b(SYNTHESIZED_WIRE_2386),
	.co(SYNTHESIZED_WIRE_2387),
	.s(SYNTHESIZED_WIRE_2279));


OneBitAdder	b2v_inst828(
	.ci(SYNTHESIZED_WIRE_2387),
	.a(SYNTHESIZED_WIRE_2388),
	.b(SYNTHESIZED_WIRE_2389),
	.co(SYNTHESIZED_WIRE_2390),
	.s(SYNTHESIZED_WIRE_2282));


OneBitAdder	b2v_inst829(
	.ci(SYNTHESIZED_WIRE_2390),
	.a(SYNTHESIZED_WIRE_2391),
	.b(SYNTHESIZED_WIRE_2392),
	.co(SYNTHESIZED_WIRE_2396),
	.s(SYNTHESIZED_WIRE_2285));


OneBitAdder	b2v_inst83(
	.ci(SYNTHESIZED_WIRE_2393),
	.a(SYNTHESIZED_WIRE_2394),
	.b(SYNTHESIZED_WIRE_2395),
	.co(SYNTHESIZED_WIRE_2425),
	.s(SYNTHESIZED_WIRE_1349));


OneBitAdder	b2v_inst830(
	.ci(SYNTHESIZED_WIRE_2396),
	.a(SYNTHESIZED_WIRE_2397),
	.b(SYNTHESIZED_WIRE_2398),
	.co(SYNTHESIZED_WIRE_2399),
	.s(SYNTHESIZED_WIRE_2288));


OneBitAdder	b2v_inst831(
	.ci(SYNTHESIZED_WIRE_2399),
	.a(SYNTHESIZED_WIRE_2400),
	.b(SYNTHESIZED_WIRE_2401),
	.co(SYNTHESIZED_WIRE_2402),
	.s(SYNTHESIZED_WIRE_2291));


OneBitAdder	b2v_inst832(
	.ci(SYNTHESIZED_WIRE_2402),
	.a(SYNTHESIZED_WIRE_2403),
	.b(SYNTHESIZED_WIRE_2404),
	.co(SYNTHESIZED_WIRE_2303),
	.s(SYNTHESIZED_WIRE_2294));


OneBitAdderHalf	b2v_inst833(
	.A(SYNTHESIZED_WIRE_2405),
	.B(SYNTHESIZED_WIRE_2406),
	.C(SYNTHESIZED_WIRE_2455),
	.S(Z_ALTERA_SYNTHESIZED[6]));


OneBitAdder	b2v_inst834(
	.ci(SYNTHESIZED_WIRE_2407),
	.a(SYNTHESIZED_WIRE_2408),
	.b(SYNTHESIZED_WIRE_2409),
	.co(SYNTHESIZED_WIRE_2410),
	.s(SYNTHESIZED_WIRE_2404));


OneBitAdder	b2v_inst835(
	.ci(SYNTHESIZED_WIRE_2410),
	.a(SYNTHESIZED_WIRE_2411),
	.b(SYNTHESIZED_WIRE_2412),
	.co(SYNTHESIZED_WIRE_2413),
	.s(SYNTHESIZED_WIRE_2305));


OneBitAdder	b2v_inst836(
	.ci(SYNTHESIZED_WIRE_2413),
	.a(SYNTHESIZED_WIRE_2414),
	.b(SYNTHESIZED_WIRE_2415),
	.co(SYNTHESIZED_WIRE_2416),
	.s(SYNTHESIZED_WIRE_2308));


OneBitAdder	b2v_inst837(
	.ci(SYNTHESIZED_WIRE_2416),
	.a(SYNTHESIZED_WIRE_2417),
	.b(SYNTHESIZED_WIRE_2418),
	.co(SYNTHESIZED_WIRE_2419),
	.s(SYNTHESIZED_WIRE_2311));


OneBitAdder	b2v_inst838(
	.ci(SYNTHESIZED_WIRE_2419),
	.a(SYNTHESIZED_WIRE_2420),
	.b(SYNTHESIZED_WIRE_2421),
	.co(SYNTHESIZED_WIRE_2422),
	.s(SYNTHESIZED_WIRE_2314));


OneBitAdder	b2v_inst839(
	.ci(SYNTHESIZED_WIRE_2422),
	.a(SYNTHESIZED_WIRE_2423),
	.b(SYNTHESIZED_WIRE_2424),
	.co(SYNTHESIZED_WIRE_2428),
	.s(SYNTHESIZED_WIRE_2317));


OneBitAdder	b2v_inst84(
	.ci(SYNTHESIZED_WIRE_2425),
	.a(SYNTHESIZED_WIRE_2426),
	.b(SYNTHESIZED_WIRE_2427),
	.co(SYNTHESIZED_WIRE_2458),
	.s(SYNTHESIZED_WIRE_1381));


OneBitAdder	b2v_inst840(
	.ci(SYNTHESIZED_WIRE_2428),
	.a(SYNTHESIZED_WIRE_2429),
	.b(SYNTHESIZED_WIRE_2430),
	.co(SYNTHESIZED_WIRE_2431),
	.s(SYNTHESIZED_WIRE_2320));


OneBitAdder	b2v_inst841(
	.ci(SYNTHESIZED_WIRE_2431),
	.a(SYNTHESIZED_WIRE_2432),
	.b(SYNTHESIZED_WIRE_2433),
	.co(SYNTHESIZED_WIRE_2434),
	.s(SYNTHESIZED_WIRE_2323));


OneBitAdder	b2v_inst842(
	.ci(SYNTHESIZED_WIRE_2434),
	.a(SYNTHESIZED_WIRE_2435),
	.b(SYNTHESIZED_WIRE_2436),
	.co(SYNTHESIZED_WIRE_2437),
	.s(SYNTHESIZED_WIRE_2326));


OneBitAdder	b2v_inst843(
	.ci(SYNTHESIZED_WIRE_2437),
	.a(SYNTHESIZED_WIRE_2438),
	.b(SYNTHESIZED_WIRE_2439),
	.co(SYNTHESIZED_WIRE_2440),
	.s(SYNTHESIZED_WIRE_2332));


OneBitAdder	b2v_inst844(
	.ci(SYNTHESIZED_WIRE_2440),
	.a(SYNTHESIZED_WIRE_2441),
	.b(SYNTHESIZED_WIRE_2442),
	.co(SYNTHESIZED_WIRE_2443),
	.s(SYNTHESIZED_WIRE_2335));


OneBitAdder	b2v_inst845(
	.ci(SYNTHESIZED_WIRE_2443),
	.a(SYNTHESIZED_WIRE_2444),
	.b(SYNTHESIZED_WIRE_2445),
	.co(SYNTHESIZED_WIRE_2446),
	.s(SYNTHESIZED_WIRE_2338));


OneBitAdder	b2v_inst846(
	.ci(SYNTHESIZED_WIRE_2446),
	.a(SYNTHESIZED_WIRE_2447),
	.b(SYNTHESIZED_WIRE_2448),
	.co(SYNTHESIZED_WIRE_2449),
	.s(SYNTHESIZED_WIRE_2341));


OneBitAdder	b2v_inst847(
	.ci(SYNTHESIZED_WIRE_2449),
	.a(SYNTHESIZED_WIRE_2450),
	.b(SYNTHESIZED_WIRE_2451),
	.co(SYNTHESIZED_WIRE_2452),
	.s(SYNTHESIZED_WIRE_2344));


OneBitAdder	b2v_inst848(
	.ci(SYNTHESIZED_WIRE_2452),
	.a(SYNTHESIZED_WIRE_2453),
	.b(SYNTHESIZED_WIRE_2454),
	.co(SYNTHESIZED_WIRE_2350),
	.s(SYNTHESIZED_WIRE_2347));


OneBitAdder	b2v_inst849(
	.ci(SYNTHESIZED_WIRE_2455),
	.a(SYNTHESIZED_WIRE_2456),
	.b(SYNTHESIZED_WIRE_2457),
	.co(SYNTHESIZED_WIRE_2461),
	.s(SYNTHESIZED_WIRE_2301));


OneBitAdder	b2v_inst85(
	.ci(SYNTHESIZED_WIRE_2458),
	.a(SYNTHESIZED_WIRE_2459),
	.b(SYNTHESIZED_WIRE_2460),
	.co(SYNTHESIZED_WIRE_2491),
	.s(SYNTHESIZED_WIRE_1414));


OneBitAdder	b2v_inst850(
	.ci(SYNTHESIZED_WIRE_2461),
	.a(SYNTHESIZED_WIRE_2462),
	.b(SYNTHESIZED_WIRE_2463),
	.co(SYNTHESIZED_WIRE_2464),
	.s(SYNTHESIZED_WIRE_2353));


OneBitAdder	b2v_inst851(
	.ci(SYNTHESIZED_WIRE_2464),
	.a(SYNTHESIZED_WIRE_2465),
	.b(SYNTHESIZED_WIRE_2466),
	.co(SYNTHESIZED_WIRE_2467),
	.s(SYNTHESIZED_WIRE_2356));


OneBitAdder	b2v_inst852(
	.ci(SYNTHESIZED_WIRE_2467),
	.a(SYNTHESIZED_WIRE_2468),
	.b(SYNTHESIZED_WIRE_2469),
	.co(SYNTHESIZED_WIRE_2470),
	.s(SYNTHESIZED_WIRE_2359));


OneBitAdder	b2v_inst853(
	.ci(SYNTHESIZED_WIRE_2470),
	.a(SYNTHESIZED_WIRE_2471),
	.b(SYNTHESIZED_WIRE_2472),
	.co(SYNTHESIZED_WIRE_2473),
	.s(SYNTHESIZED_WIRE_2365));


OneBitAdder	b2v_inst854(
	.ci(SYNTHESIZED_WIRE_2473),
	.a(SYNTHESIZED_WIRE_2474),
	.b(SYNTHESIZED_WIRE_2475),
	.co(SYNTHESIZED_WIRE_2476),
	.s(SYNTHESIZED_WIRE_2368));


OneBitAdder	b2v_inst855(
	.ci(SYNTHESIZED_WIRE_2476),
	.a(SYNTHESIZED_WIRE_2477),
	.b(SYNTHESIZED_WIRE_2478),
	.co(SYNTHESIZED_WIRE_2479),
	.s(SYNTHESIZED_WIRE_2371));


OneBitAdder	b2v_inst856(
	.ci(SYNTHESIZED_WIRE_2479),
	.a(SYNTHESIZED_WIRE_2480),
	.b(SYNTHESIZED_WIRE_2481),
	.co(SYNTHESIZED_WIRE_2482),
	.s(SYNTHESIZED_WIRE_2374));


OneBitAdder	b2v_inst857(
	.ci(SYNTHESIZED_WIRE_2482),
	.a(SYNTHESIZED_WIRE_2483),
	.b(SYNTHESIZED_WIRE_2484),
	.co(SYNTHESIZED_WIRE_2485),
	.s(SYNTHESIZED_WIRE_2377));


OneBitAdder	b2v_inst858(
	.ci(SYNTHESIZED_WIRE_2485),
	.a(SYNTHESIZED_WIRE_2486),
	.b(SYNTHESIZED_WIRE_2487),
	.co(SYNTHESIZED_WIRE_2488),
	.s(SYNTHESIZED_WIRE_2380));


OneBitAdder	b2v_inst859(
	.ci(SYNTHESIZED_WIRE_2488),
	.a(SYNTHESIZED_WIRE_2489),
	.b(SYNTHESIZED_WIRE_2490),
	.co(SYNTHESIZED_WIRE_2494),
	.s(SYNTHESIZED_WIRE_2383));


OneBitAdder	b2v_inst86(
	.ci(SYNTHESIZED_WIRE_2491),
	.a(SYNTHESIZED_WIRE_2492),
	.b(SYNTHESIZED_WIRE_2493),
	.co(SYNTHESIZED_WIRE_2523),
	.s(SYNTHESIZED_WIRE_1447));


OneBitAdder	b2v_inst860(
	.ci(SYNTHESIZED_WIRE_2494),
	.a(SYNTHESIZED_WIRE_2495),
	.b(SYNTHESIZED_WIRE_2496),
	.co(SYNTHESIZED_WIRE_2497),
	.s(SYNTHESIZED_WIRE_2386));


OneBitAdder	b2v_inst861(
	.ci(SYNTHESIZED_WIRE_2497),
	.a(SYNTHESIZED_WIRE_2498),
	.b(SYNTHESIZED_WIRE_2499),
	.co(SYNTHESIZED_WIRE_2500),
	.s(SYNTHESIZED_WIRE_2389));


OneBitAdder	b2v_inst862(
	.ci(SYNTHESIZED_WIRE_2500),
	.a(SYNTHESIZED_WIRE_2501),
	.b(SYNTHESIZED_WIRE_2502),
	.co(SYNTHESIZED_WIRE_2503),
	.s(SYNTHESIZED_WIRE_2392));


OneBitAdder	b2v_inst863(
	.ci(SYNTHESIZED_WIRE_2503),
	.a(SYNTHESIZED_WIRE_2504),
	.b(SYNTHESIZED_WIRE_2505),
	.co(SYNTHESIZED_WIRE_2506),
	.s(SYNTHESIZED_WIRE_2398));


OneBitAdder	b2v_inst864(
	.ci(SYNTHESIZED_WIRE_2506),
	.a(SYNTHESIZED_WIRE_2507),
	.b(SYNTHESIZED_WIRE_2508),
	.co(SYNTHESIZED_WIRE_2407),
	.s(SYNTHESIZED_WIRE_2401));


OneBitAdderHalf	b2v_inst865(
	.A(SYNTHESIZED_WIRE_2509),
	.B(SYNTHESIZED_WIRE_2510),
	.C(SYNTHESIZED_WIRE_2562),
	.S(Z_ALTERA_SYNTHESIZED[5]));


OneBitAdder	b2v_inst866(
	.ci(SYNTHESIZED_WIRE_2511),
	.a(SYNTHESIZED_WIRE_2512),
	.b(SYNTHESIZED_WIRE_2513),
	.co(SYNTHESIZED_WIRE_2514),
	.s(SYNTHESIZED_WIRE_2508));


OneBitAdder	b2v_inst867(
	.ci(SYNTHESIZED_WIRE_2514),
	.a(SYNTHESIZED_WIRE_2515),
	.b(SYNTHESIZED_WIRE_2516),
	.co(SYNTHESIZED_WIRE_2517),
	.s(SYNTHESIZED_WIRE_2409));


OneBitAdder	b2v_inst868(
	.ci(SYNTHESIZED_WIRE_2517),
	.a(SYNTHESIZED_WIRE_2518),
	.b(SYNTHESIZED_WIRE_2519),
	.co(SYNTHESIZED_WIRE_2520),
	.s(SYNTHESIZED_WIRE_2412));


OneBitAdder	b2v_inst869(
	.ci(SYNTHESIZED_WIRE_2520),
	.a(SYNTHESIZED_WIRE_2521),
	.b(SYNTHESIZED_WIRE_2522),
	.co(SYNTHESIZED_WIRE_2526),
	.s(SYNTHESIZED_WIRE_2415));


OneBitAdder	b2v_inst87(
	.ci(SYNTHESIZED_WIRE_2523),
	.a(SYNTHESIZED_WIRE_2524),
	.b(SYNTHESIZED_WIRE_2525),
	.co(SYNTHESIZED_WIRE_2556),
	.s(SYNTHESIZED_WIRE_1479));


OneBitAdder	b2v_inst870(
	.ci(SYNTHESIZED_WIRE_2526),
	.a(SYNTHESIZED_WIRE_2527),
	.b(SYNTHESIZED_WIRE_2528),
	.co(SYNTHESIZED_WIRE_2529),
	.s(SYNTHESIZED_WIRE_2418));


OneBitAdder	b2v_inst871(
	.ci(SYNTHESIZED_WIRE_2529),
	.a(SYNTHESIZED_WIRE_2530),
	.b(SYNTHESIZED_WIRE_2531),
	.co(SYNTHESIZED_WIRE_2532),
	.s(SYNTHESIZED_WIRE_2421));


OneBitAdder	b2v_inst872(
	.ci(SYNTHESIZED_WIRE_2532),
	.a(SYNTHESIZED_WIRE_2533),
	.b(SYNTHESIZED_WIRE_2534),
	.co(SYNTHESIZED_WIRE_2535),
	.s(SYNTHESIZED_WIRE_2424));


OneBitAdder	b2v_inst873(
	.ci(SYNTHESIZED_WIRE_2535),
	.a(SYNTHESIZED_WIRE_2536),
	.b(SYNTHESIZED_WIRE_2537),
	.co(SYNTHESIZED_WIRE_2538),
	.s(SYNTHESIZED_WIRE_2430));


OneBitAdder	b2v_inst874(
	.ci(SYNTHESIZED_WIRE_2538),
	.a(SYNTHESIZED_WIRE_2539),
	.b(SYNTHESIZED_WIRE_2540),
	.co(SYNTHESIZED_WIRE_2541),
	.s(SYNTHESIZED_WIRE_2433));


OneBitAdder	b2v_inst875(
	.ci(SYNTHESIZED_WIRE_2541),
	.a(SYNTHESIZED_WIRE_2542),
	.b(SYNTHESIZED_WIRE_2543),
	.co(SYNTHESIZED_WIRE_2544),
	.s(SYNTHESIZED_WIRE_2436));


OneBitAdder	b2v_inst876(
	.ci(SYNTHESIZED_WIRE_2544),
	.a(SYNTHESIZED_WIRE_2545),
	.b(SYNTHESIZED_WIRE_2546),
	.co(SYNTHESIZED_WIRE_2547),
	.s(SYNTHESIZED_WIRE_2439));


OneBitAdder	b2v_inst877(
	.ci(SYNTHESIZED_WIRE_2547),
	.a(SYNTHESIZED_WIRE_2548),
	.b(SYNTHESIZED_WIRE_2549),
	.co(SYNTHESIZED_WIRE_2550),
	.s(SYNTHESIZED_WIRE_2442));


OneBitAdder	b2v_inst878(
	.ci(SYNTHESIZED_WIRE_2550),
	.a(SYNTHESIZED_WIRE_2551),
	.b(SYNTHESIZED_WIRE_2552),
	.co(SYNTHESIZED_WIRE_2553),
	.s(SYNTHESIZED_WIRE_2445));


OneBitAdder	b2v_inst879(
	.ci(SYNTHESIZED_WIRE_2553),
	.a(SYNTHESIZED_WIRE_2554),
	.b(SYNTHESIZED_WIRE_2555),
	.co(SYNTHESIZED_WIRE_2559),
	.s(SYNTHESIZED_WIRE_2448));


OneBitAdder	b2v_inst88(
	.ci(SYNTHESIZED_WIRE_2556),
	.a(SYNTHESIZED_WIRE_2557),
	.b(SYNTHESIZED_WIRE_2558),
	.co(SYNTHESIZED_WIRE_2589),
	.s(SYNTHESIZED_WIRE_1512));


OneBitAdder	b2v_inst880(
	.ci(SYNTHESIZED_WIRE_2559),
	.a(SYNTHESIZED_WIRE_2560),
	.b(SYNTHESIZED_WIRE_2561),
	.co(SYNTHESIZED_WIRE_2454),
	.s(SYNTHESIZED_WIRE_2451));


OneBitAdder	b2v_inst881(
	.ci(SYNTHESIZED_WIRE_2562),
	.a(SYNTHESIZED_WIRE_2563),
	.b(SYNTHESIZED_WIRE_2564),
	.co(SYNTHESIZED_WIRE_2565),
	.s(SYNTHESIZED_WIRE_2405));


OneBitAdder	b2v_inst882(
	.ci(SYNTHESIZED_WIRE_2565),
	.a(SYNTHESIZED_WIRE_2566),
	.b(SYNTHESIZED_WIRE_2567),
	.co(SYNTHESIZED_WIRE_2568),
	.s(SYNTHESIZED_WIRE_2457));


OneBitAdder	b2v_inst883(
	.ci(SYNTHESIZED_WIRE_2568),
	.a(SYNTHESIZED_WIRE_2569),
	.b(SYNTHESIZED_WIRE_2570),
	.co(SYNTHESIZED_WIRE_2571),
	.s(SYNTHESIZED_WIRE_2463));


OneBitAdder	b2v_inst884(
	.ci(SYNTHESIZED_WIRE_2571),
	.a(SYNTHESIZED_WIRE_2572),
	.b(SYNTHESIZED_WIRE_2573),
	.co(SYNTHESIZED_WIRE_2574),
	.s(SYNTHESIZED_WIRE_2466));


OneBitAdder	b2v_inst885(
	.ci(SYNTHESIZED_WIRE_2574),
	.a(SYNTHESIZED_WIRE_2575),
	.b(SYNTHESIZED_WIRE_2576),
	.co(SYNTHESIZED_WIRE_2577),
	.s(SYNTHESIZED_WIRE_2469));


OneBitAdder	b2v_inst886(
	.ci(SYNTHESIZED_WIRE_2577),
	.a(SYNTHESIZED_WIRE_2578),
	.b(SYNTHESIZED_WIRE_2579),
	.co(SYNTHESIZED_WIRE_2580),
	.s(SYNTHESIZED_WIRE_2472));


OneBitAdder	b2v_inst887(
	.ci(SYNTHESIZED_WIRE_2580),
	.a(SYNTHESIZED_WIRE_2581),
	.b(SYNTHESIZED_WIRE_2582),
	.co(SYNTHESIZED_WIRE_2583),
	.s(SYNTHESIZED_WIRE_2475));


OneBitAdder	b2v_inst888(
	.ci(SYNTHESIZED_WIRE_2583),
	.a(SYNTHESIZED_WIRE_2584),
	.b(SYNTHESIZED_WIRE_2585),
	.co(SYNTHESIZED_WIRE_2586),
	.s(SYNTHESIZED_WIRE_2478));


OneBitAdder	b2v_inst889(
	.ci(SYNTHESIZED_WIRE_2586),
	.a(SYNTHESIZED_WIRE_2587),
	.b(SYNTHESIZED_WIRE_2588),
	.co(SYNTHESIZED_WIRE_2592),
	.s(SYNTHESIZED_WIRE_2481));


OneBitAdder	b2v_inst89(
	.ci(SYNTHESIZED_WIRE_2589),
	.a(SYNTHESIZED_WIRE_2590),
	.b(SYNTHESIZED_WIRE_2591),
	.co(SYNTHESIZED_WIRE_2621),
	.s(SYNTHESIZED_WIRE_1545));


OneBitAdder	b2v_inst890(
	.ci(SYNTHESIZED_WIRE_2592),
	.a(SYNTHESIZED_WIRE_2593),
	.b(SYNTHESIZED_WIRE_2594),
	.co(SYNTHESIZED_WIRE_2595),
	.s(SYNTHESIZED_WIRE_2484));


OneBitAdder	b2v_inst891(
	.ci(SYNTHESIZED_WIRE_2595),
	.a(SYNTHESIZED_WIRE_2596),
	.b(SYNTHESIZED_WIRE_2597),
	.co(SYNTHESIZED_WIRE_2598),
	.s(SYNTHESIZED_WIRE_2487));


OneBitAdder	b2v_inst892(
	.ci(SYNTHESIZED_WIRE_2598),
	.a(SYNTHESIZED_WIRE_2599),
	.b(SYNTHESIZED_WIRE_2600),
	.co(SYNTHESIZED_WIRE_2601),
	.s(SYNTHESIZED_WIRE_2490));


OneBitAdder	b2v_inst893(
	.ci(SYNTHESIZED_WIRE_2601),
	.a(SYNTHESIZED_WIRE_2602),
	.b(SYNTHESIZED_WIRE_2603),
	.co(SYNTHESIZED_WIRE_2604),
	.s(SYNTHESIZED_WIRE_2496));


OneBitAdder	b2v_inst894(
	.ci(SYNTHESIZED_WIRE_2604),
	.a(SYNTHESIZED_WIRE_2605),
	.b(SYNTHESIZED_WIRE_2606),
	.co(SYNTHESIZED_WIRE_2607),
	.s(SYNTHESIZED_WIRE_2499));


OneBitAdder	b2v_inst895(
	.ci(SYNTHESIZED_WIRE_2607),
	.a(SYNTHESIZED_WIRE_2608),
	.b(SYNTHESIZED_WIRE_2609),
	.co(SYNTHESIZED_WIRE_2610),
	.s(SYNTHESIZED_WIRE_2502));


OneBitAdder	b2v_inst896(
	.ci(SYNTHESIZED_WIRE_2610),
	.a(SYNTHESIZED_WIRE_2611),
	.b(SYNTHESIZED_WIRE_2612),
	.co(SYNTHESIZED_WIRE_2511),
	.s(SYNTHESIZED_WIRE_2505));


OneBitAdderHalf	b2v_inst897(
	.A(SYNTHESIZED_WIRE_2613),
	.B(SYNTHESIZED_WIRE_2614),
	.C(SYNTHESIZED_WIRE_2666),
	.S(Z_ALTERA_SYNTHESIZED[4]));


OneBitAdder	b2v_inst898(
	.ci(SYNTHESIZED_WIRE_2615),
	.a(SYNTHESIZED_WIRE_2616),
	.b(SYNTHESIZED_WIRE_2617),
	.co(SYNTHESIZED_WIRE_2618),
	.s(SYNTHESIZED_WIRE_2612));


OneBitAdder	b2v_inst899(
	.ci(SYNTHESIZED_WIRE_2618),
	.a(SYNTHESIZED_WIRE_2619),
	.b(SYNTHESIZED_WIRE_2620),
	.co(SYNTHESIZED_WIRE_2624),
	.s(SYNTHESIZED_WIRE_2513));


OneBitAdder	b2v_inst90(
	.ci(SYNTHESIZED_WIRE_2621),
	.a(SYNTHESIZED_WIRE_2622),
	.b(SYNTHESIZED_WIRE_2623),
	.co(SYNTHESIZED_WIRE_2654),
	.s(SYNTHESIZED_WIRE_1577));


OneBitAdder	b2v_inst900(
	.ci(SYNTHESIZED_WIRE_2624),
	.a(SYNTHESIZED_WIRE_2625),
	.b(SYNTHESIZED_WIRE_2626),
	.co(SYNTHESIZED_WIRE_2627),
	.s(SYNTHESIZED_WIRE_2516));


OneBitAdder	b2v_inst901(
	.ci(SYNTHESIZED_WIRE_2627),
	.a(SYNTHESIZED_WIRE_2628),
	.b(SYNTHESIZED_WIRE_2629),
	.co(SYNTHESIZED_WIRE_2630),
	.s(SYNTHESIZED_WIRE_2519));


OneBitAdder	b2v_inst902(
	.ci(SYNTHESIZED_WIRE_2630),
	.a(SYNTHESIZED_WIRE_2631),
	.b(SYNTHESIZED_WIRE_2632),
	.co(SYNTHESIZED_WIRE_2633),
	.s(SYNTHESIZED_WIRE_2522));


OneBitAdder	b2v_inst903(
	.ci(SYNTHESIZED_WIRE_2633),
	.a(SYNTHESIZED_WIRE_2634),
	.b(SYNTHESIZED_WIRE_2635),
	.co(SYNTHESIZED_WIRE_2636),
	.s(SYNTHESIZED_WIRE_2528));


OneBitAdder	b2v_inst904(
	.ci(SYNTHESIZED_WIRE_2636),
	.a(SYNTHESIZED_WIRE_2637),
	.b(SYNTHESIZED_WIRE_2638),
	.co(SYNTHESIZED_WIRE_2639),
	.s(SYNTHESIZED_WIRE_2531));


OneBitAdder	b2v_inst905(
	.ci(SYNTHESIZED_WIRE_2639),
	.a(SYNTHESIZED_WIRE_2640),
	.b(SYNTHESIZED_WIRE_2641),
	.co(SYNTHESIZED_WIRE_2642),
	.s(SYNTHESIZED_WIRE_2534));


OneBitAdder	b2v_inst906(
	.ci(SYNTHESIZED_WIRE_2642),
	.a(SYNTHESIZED_WIRE_2643),
	.b(SYNTHESIZED_WIRE_2644),
	.co(SYNTHESIZED_WIRE_2645),
	.s(SYNTHESIZED_WIRE_2537));


OneBitAdder	b2v_inst907(
	.ci(SYNTHESIZED_WIRE_2645),
	.a(SYNTHESIZED_WIRE_2646),
	.b(SYNTHESIZED_WIRE_2647),
	.co(SYNTHESIZED_WIRE_2648),
	.s(SYNTHESIZED_WIRE_2540));


OneBitAdder	b2v_inst908(
	.ci(SYNTHESIZED_WIRE_2648),
	.a(SYNTHESIZED_WIRE_2649),
	.b(SYNTHESIZED_WIRE_2650),
	.co(SYNTHESIZED_WIRE_2651),
	.s(SYNTHESIZED_WIRE_2543));


OneBitAdder	b2v_inst909(
	.ci(SYNTHESIZED_WIRE_2651),
	.a(SYNTHESIZED_WIRE_2652),
	.b(SYNTHESIZED_WIRE_2653),
	.co(SYNTHESIZED_WIRE_2657),
	.s(SYNTHESIZED_WIRE_2546));


OneBitAdder	b2v_inst91(
	.ci(SYNTHESIZED_WIRE_2654),
	.a(SYNTHESIZED_WIRE_2655),
	.b(SYNTHESIZED_WIRE_2656),
	.co(SYNTHESIZED_WIRE_2687),
	.s(SYNTHESIZED_WIRE_1610));


OneBitAdder	b2v_inst910(
	.ci(SYNTHESIZED_WIRE_2657),
	.a(SYNTHESIZED_WIRE_2658),
	.b(SYNTHESIZED_WIRE_2659),
	.co(SYNTHESIZED_WIRE_2660),
	.s(SYNTHESIZED_WIRE_2549));


OneBitAdder	b2v_inst911(
	.ci(SYNTHESIZED_WIRE_2660),
	.a(SYNTHESIZED_WIRE_2661),
	.b(SYNTHESIZED_WIRE_2662),
	.co(SYNTHESIZED_WIRE_2663),
	.s(SYNTHESIZED_WIRE_2552));


OneBitAdder	b2v_inst912(
	.ci(SYNTHESIZED_WIRE_2663),
	.a(SYNTHESIZED_WIRE_2664),
	.b(SYNTHESIZED_WIRE_2665),
	.co(SYNTHESIZED_WIRE_2561),
	.s(SYNTHESIZED_WIRE_2555));


OneBitAdder	b2v_inst913(
	.ci(SYNTHESIZED_WIRE_2666),
	.a(SYNTHESIZED_WIRE_2667),
	.b(SYNTHESIZED_WIRE_2668),
	.co(SYNTHESIZED_WIRE_2669),
	.s(SYNTHESIZED_WIRE_2509));


OneBitAdder	b2v_inst914(
	.ci(SYNTHESIZED_WIRE_2669),
	.a(SYNTHESIZED_WIRE_2670),
	.b(SYNTHESIZED_WIRE_2671),
	.co(SYNTHESIZED_WIRE_2672),
	.s(SYNTHESIZED_WIRE_2564));


OneBitAdder	b2v_inst915(
	.ci(SYNTHESIZED_WIRE_2672),
	.a(SYNTHESIZED_WIRE_2673),
	.b(SYNTHESIZED_WIRE_2674),
	.co(SYNTHESIZED_WIRE_2675),
	.s(SYNTHESIZED_WIRE_2567));


OneBitAdder	b2v_inst916(
	.ci(SYNTHESIZED_WIRE_2675),
	.a(SYNTHESIZED_WIRE_2676),
	.b(SYNTHESIZED_WIRE_2677),
	.co(SYNTHESIZED_WIRE_2678),
	.s(SYNTHESIZED_WIRE_2570));


OneBitAdder	b2v_inst917(
	.ci(SYNTHESIZED_WIRE_2678),
	.a(SYNTHESIZED_WIRE_2679),
	.b(SYNTHESIZED_WIRE_2680),
	.co(SYNTHESIZED_WIRE_2681),
	.s(SYNTHESIZED_WIRE_2573));


OneBitAdder	b2v_inst918(
	.ci(SYNTHESIZED_WIRE_2681),
	.a(SYNTHESIZED_WIRE_2682),
	.b(SYNTHESIZED_WIRE_2683),
	.co(SYNTHESIZED_WIRE_2684),
	.s(SYNTHESIZED_WIRE_2576));


OneBitAdder	b2v_inst919(
	.ci(SYNTHESIZED_WIRE_2684),
	.a(SYNTHESIZED_WIRE_2685),
	.b(SYNTHESIZED_WIRE_2686),
	.co(SYNTHESIZED_WIRE_2690),
	.s(SYNTHESIZED_WIRE_2579));


OneBitAdder	b2v_inst92(
	.ci(SYNTHESIZED_WIRE_2687),
	.a(SYNTHESIZED_WIRE_2688),
	.b(SYNTHESIZED_WIRE_2689),
	.co(SYNTHESIZED_WIRE_2719),
	.s(SYNTHESIZED_WIRE_1643));


OneBitAdder	b2v_inst920(
	.ci(SYNTHESIZED_WIRE_2690),
	.a(SYNTHESIZED_WIRE_2691),
	.b(SYNTHESIZED_WIRE_2692),
	.co(SYNTHESIZED_WIRE_2693),
	.s(SYNTHESIZED_WIRE_2582));


OneBitAdder	b2v_inst921(
	.ci(SYNTHESIZED_WIRE_2693),
	.a(SYNTHESIZED_WIRE_2694),
	.b(SYNTHESIZED_WIRE_2695),
	.co(SYNTHESIZED_WIRE_2696),
	.s(SYNTHESIZED_WIRE_2585));


OneBitAdder	b2v_inst922(
	.ci(SYNTHESIZED_WIRE_2696),
	.a(SYNTHESIZED_WIRE_2697),
	.b(SYNTHESIZED_WIRE_2698),
	.co(SYNTHESIZED_WIRE_2699),
	.s(SYNTHESIZED_WIRE_2588));


OneBitAdder	b2v_inst923(
	.ci(SYNTHESIZED_WIRE_2699),
	.a(SYNTHESIZED_WIRE_2700),
	.b(SYNTHESIZED_WIRE_2701),
	.co(SYNTHESIZED_WIRE_2702),
	.s(SYNTHESIZED_WIRE_2594));


OneBitAdder	b2v_inst924(
	.ci(SYNTHESIZED_WIRE_2702),
	.a(SYNTHESIZED_WIRE_2703),
	.b(SYNTHESIZED_WIRE_2704),
	.co(SYNTHESIZED_WIRE_2705),
	.s(SYNTHESIZED_WIRE_2597));


OneBitAdder	b2v_inst925(
	.ci(SYNTHESIZED_WIRE_2705),
	.a(SYNTHESIZED_WIRE_2706),
	.b(SYNTHESIZED_WIRE_2707),
	.co(SYNTHESIZED_WIRE_2708),
	.s(SYNTHESIZED_WIRE_2600));


OneBitAdder	b2v_inst926(
	.ci(SYNTHESIZED_WIRE_2708),
	.a(SYNTHESIZED_WIRE_2709),
	.b(SYNTHESIZED_WIRE_2710),
	.co(SYNTHESIZED_WIRE_2711),
	.s(SYNTHESIZED_WIRE_2603));


OneBitAdder	b2v_inst927(
	.ci(SYNTHESIZED_WIRE_2711),
	.a(SYNTHESIZED_WIRE_2712),
	.b(SYNTHESIZED_WIRE_2713),
	.co(SYNTHESIZED_WIRE_2714),
	.s(SYNTHESIZED_WIRE_2606));


OneBitAdder	b2v_inst928(
	.ci(SYNTHESIZED_WIRE_2714),
	.a(SYNTHESIZED_WIRE_2715),
	.b(SYNTHESIZED_WIRE_2716),
	.co(SYNTHESIZED_WIRE_2615),
	.s(SYNTHESIZED_WIRE_2609));


OneBitAdderHalf	b2v_inst929(
	.A(SYNTHESIZED_WIRE_2717),
	.B(SYNTHESIZED_WIRE_2718),
	.C(SYNTHESIZED_WIRE_2770),
	.S(Z_ALTERA_SYNTHESIZED[3]));


OneBitAdder	b2v_inst93(
	.ci(SYNTHESIZED_WIRE_2719),
	.a(SYNTHESIZED_WIRE_2720),
	.b(SYNTHESIZED_WIRE_2721),
	.co(SYNTHESIZED_WIRE_2752),
	.s(SYNTHESIZED_WIRE_1675));


OneBitAdder	b2v_inst930(
	.ci(SYNTHESIZED_WIRE_2722),
	.a(SYNTHESIZED_WIRE_2723),
	.b(SYNTHESIZED_WIRE_2724),
	.co(SYNTHESIZED_WIRE_2725),
	.s(SYNTHESIZED_WIRE_2716));


OneBitAdder	b2v_inst931(
	.ci(SYNTHESIZED_WIRE_2725),
	.a(SYNTHESIZED_WIRE_2726),
	.b(SYNTHESIZED_WIRE_2727),
	.co(SYNTHESIZED_WIRE_2728),
	.s(SYNTHESIZED_WIRE_2617));


OneBitAdder	b2v_inst932(
	.ci(SYNTHESIZED_WIRE_2728),
	.a(SYNTHESIZED_WIRE_2729),
	.b(SYNTHESIZED_WIRE_2730),
	.co(SYNTHESIZED_WIRE_2731),
	.s(SYNTHESIZED_WIRE_2620));


OneBitAdder	b2v_inst933(
	.ci(SYNTHESIZED_WIRE_2731),
	.a(SYNTHESIZED_WIRE_2732),
	.b(SYNTHESIZED_WIRE_2733),
	.co(SYNTHESIZED_WIRE_2734),
	.s(SYNTHESIZED_WIRE_2626));


OneBitAdder	b2v_inst934(
	.ci(SYNTHESIZED_WIRE_2734),
	.a(SYNTHESIZED_WIRE_2735),
	.b(SYNTHESIZED_WIRE_2736),
	.co(SYNTHESIZED_WIRE_2737),
	.s(SYNTHESIZED_WIRE_2629));


OneBitAdder	b2v_inst935(
	.ci(SYNTHESIZED_WIRE_2737),
	.a(SYNTHESIZED_WIRE_2738),
	.b(SYNTHESIZED_WIRE_2739),
	.co(SYNTHESIZED_WIRE_2740),
	.s(SYNTHESIZED_WIRE_2632));


OneBitAdder	b2v_inst936(
	.ci(SYNTHESIZED_WIRE_2740),
	.a(SYNTHESIZED_WIRE_2741),
	.b(SYNTHESIZED_WIRE_2742),
	.co(SYNTHESIZED_WIRE_2743),
	.s(SYNTHESIZED_WIRE_2635));


OneBitAdder	b2v_inst937(
	.ci(SYNTHESIZED_WIRE_2743),
	.a(SYNTHESIZED_WIRE_2744),
	.b(SYNTHESIZED_WIRE_2745),
	.co(SYNTHESIZED_WIRE_2746),
	.s(SYNTHESIZED_WIRE_2638));


OneBitAdder	b2v_inst938(
	.ci(SYNTHESIZED_WIRE_2746),
	.a(SYNTHESIZED_WIRE_2747),
	.b(SYNTHESIZED_WIRE_2748),
	.co(SYNTHESIZED_WIRE_2749),
	.s(SYNTHESIZED_WIRE_2641));


OneBitAdder	b2v_inst939(
	.ci(SYNTHESIZED_WIRE_2749),
	.a(SYNTHESIZED_WIRE_2750),
	.b(SYNTHESIZED_WIRE_2751),
	.co(SYNTHESIZED_WIRE_2755),
	.s(SYNTHESIZED_WIRE_2644));


OneBitAdder	b2v_inst94(
	.ci(SYNTHESIZED_WIRE_2752),
	.a(SYNTHESIZED_WIRE_2753),
	.b(SYNTHESIZED_WIRE_2754),
	.co(SYNTHESIZED_WIRE_2785),
	.s(SYNTHESIZED_WIRE_1708));


OneBitAdder	b2v_inst940(
	.ci(SYNTHESIZED_WIRE_2755),
	.a(SYNTHESIZED_WIRE_2756),
	.b(SYNTHESIZED_WIRE_2757),
	.co(SYNTHESIZED_WIRE_2758),
	.s(SYNTHESIZED_WIRE_2647));


OneBitAdder	b2v_inst941(
	.ci(SYNTHESIZED_WIRE_2758),
	.a(SYNTHESIZED_WIRE_2759),
	.b(SYNTHESIZED_WIRE_2760),
	.co(SYNTHESIZED_WIRE_2761),
	.s(SYNTHESIZED_WIRE_2650));


OneBitAdder	b2v_inst942(
	.ci(SYNTHESIZED_WIRE_2761),
	.a(SYNTHESIZED_WIRE_2762),
	.b(SYNTHESIZED_WIRE_2763),
	.co(SYNTHESIZED_WIRE_2764),
	.s(SYNTHESIZED_WIRE_2653));


OneBitAdder	b2v_inst943(
	.ci(SYNTHESIZED_WIRE_2764),
	.a(SYNTHESIZED_WIRE_2765),
	.b(SYNTHESIZED_WIRE_2766),
	.co(SYNTHESIZED_WIRE_2767),
	.s(SYNTHESIZED_WIRE_2659));


OneBitAdder	b2v_inst944(
	.ci(SYNTHESIZED_WIRE_2767),
	.a(SYNTHESIZED_WIRE_2768),
	.b(SYNTHESIZED_WIRE_2769),
	.co(SYNTHESIZED_WIRE_2665),
	.s(SYNTHESIZED_WIRE_2662));


OneBitAdder	b2v_inst945(
	.ci(SYNTHESIZED_WIRE_2770),
	.a(SYNTHESIZED_WIRE_2771),
	.b(SYNTHESIZED_WIRE_2772),
	.co(SYNTHESIZED_WIRE_2773),
	.s(SYNTHESIZED_WIRE_2613));


OneBitAdder	b2v_inst946(
	.ci(SYNTHESIZED_WIRE_2773),
	.a(SYNTHESIZED_WIRE_2774),
	.b(SYNTHESIZED_WIRE_2775),
	.co(SYNTHESIZED_WIRE_2776),
	.s(SYNTHESIZED_WIRE_2668));


OneBitAdder	b2v_inst947(
	.ci(SYNTHESIZED_WIRE_2776),
	.a(SYNTHESIZED_WIRE_2777),
	.b(SYNTHESIZED_WIRE_2778),
	.co(SYNTHESIZED_WIRE_2779),
	.s(SYNTHESIZED_WIRE_2671));


OneBitAdder	b2v_inst948(
	.ci(SYNTHESIZED_WIRE_2779),
	.a(SYNTHESIZED_WIRE_2780),
	.b(SYNTHESIZED_WIRE_2781),
	.co(SYNTHESIZED_WIRE_2782),
	.s(SYNTHESIZED_WIRE_2674));


OneBitAdder	b2v_inst949(
	.ci(SYNTHESIZED_WIRE_2782),
	.a(SYNTHESIZED_WIRE_2783),
	.b(SYNTHESIZED_WIRE_2784),
	.co(SYNTHESIZED_WIRE_2788),
	.s(SYNTHESIZED_WIRE_2677));


OneBitAdder	b2v_inst95(
	.ci(SYNTHESIZED_WIRE_2785),
	.a(SYNTHESIZED_WIRE_2786),
	.b(SYNTHESIZED_WIRE_2787),
	.co(SYNTHESIZED_WIRE_2818),
	.s(SYNTHESIZED_WIRE_1741));


OneBitAdder	b2v_inst950(
	.ci(SYNTHESIZED_WIRE_2788),
	.a(SYNTHESIZED_WIRE_2789),
	.b(SYNTHESIZED_WIRE_2790),
	.co(SYNTHESIZED_WIRE_2791),
	.s(SYNTHESIZED_WIRE_2680));


OneBitAdder	b2v_inst951(
	.ci(SYNTHESIZED_WIRE_2791),
	.a(SYNTHESIZED_WIRE_2792),
	.b(SYNTHESIZED_WIRE_2793),
	.co(SYNTHESIZED_WIRE_2794),
	.s(SYNTHESIZED_WIRE_2683));


OneBitAdder	b2v_inst952(
	.ci(SYNTHESIZED_WIRE_2794),
	.a(SYNTHESIZED_WIRE_2795),
	.b(SYNTHESIZED_WIRE_2796),
	.co(SYNTHESIZED_WIRE_2797),
	.s(SYNTHESIZED_WIRE_2686));


OneBitAdder	b2v_inst953(
	.ci(SYNTHESIZED_WIRE_2797),
	.a(SYNTHESIZED_WIRE_2798),
	.b(SYNTHESIZED_WIRE_2799),
	.co(SYNTHESIZED_WIRE_2800),
	.s(SYNTHESIZED_WIRE_2692));


OneBitAdder	b2v_inst954(
	.ci(SYNTHESIZED_WIRE_2800),
	.a(SYNTHESIZED_WIRE_2801),
	.b(SYNTHESIZED_WIRE_2802),
	.co(SYNTHESIZED_WIRE_2803),
	.s(SYNTHESIZED_WIRE_2695));


OneBitAdder	b2v_inst955(
	.ci(SYNTHESIZED_WIRE_2803),
	.a(SYNTHESIZED_WIRE_2804),
	.b(SYNTHESIZED_WIRE_2805),
	.co(SYNTHESIZED_WIRE_2806),
	.s(SYNTHESIZED_WIRE_2698));


OneBitAdder	b2v_inst956(
	.ci(SYNTHESIZED_WIRE_2806),
	.a(SYNTHESIZED_WIRE_2807),
	.b(SYNTHESIZED_WIRE_2808),
	.co(SYNTHESIZED_WIRE_2809),
	.s(SYNTHESIZED_WIRE_2701));


OneBitAdder	b2v_inst957(
	.ci(SYNTHESIZED_WIRE_2809),
	.a(SYNTHESIZED_WIRE_2810),
	.b(SYNTHESIZED_WIRE_2811),
	.co(SYNTHESIZED_WIRE_2812),
	.s(SYNTHESIZED_WIRE_2704));


OneBitAdder	b2v_inst958(
	.ci(SYNTHESIZED_WIRE_2812),
	.a(SYNTHESIZED_WIRE_2813),
	.b(SYNTHESIZED_WIRE_2814),
	.co(SYNTHESIZED_WIRE_2815),
	.s(SYNTHESIZED_WIRE_2707));


OneBitAdder	b2v_inst959(
	.ci(SYNTHESIZED_WIRE_2815),
	.a(SYNTHESIZED_WIRE_2816),
	.b(SYNTHESIZED_WIRE_2817),
	.co(SYNTHESIZED_WIRE_2821),
	.s(SYNTHESIZED_WIRE_2710));


OneBitAdder	b2v_inst96(
	.ci(SYNTHESIZED_WIRE_2818),
	.a(SYNTHESIZED_WIRE_2819),
	.b(SYNTHESIZED_WIRE_2820),
	.co(SYNTHESIZED_WIRE_1837),
	.s(SYNTHESIZED_WIRE_1774));


OneBitAdder	b2v_inst960(
	.ci(SYNTHESIZED_WIRE_2821),
	.a(SYNTHESIZED_WIRE_2822),
	.b(SYNTHESIZED_WIRE_2823),
	.co(SYNTHESIZED_WIRE_2722),
	.s(SYNTHESIZED_WIRE_2713));


OneBitAdderHalf	b2v_inst961(
	.A(SYNTHESIZED_WIRE_2824),
	.B(SYNTHESIZED_WIRE_2825),
	.C(SYNTHESIZED_WIRE_2873),
	.S(Z_ALTERA_SYNTHESIZED[2]));


OneBitAdder	b2v_inst962(
	.ci(SYNTHESIZED_WIRE_2826),
	.a(SYNTHESIZED_WIRE_2827),
	.b(SYNTHESIZED_WIRE_2828),
	.co(SYNTHESIZED_WIRE_2829),
	.s(SYNTHESIZED_WIRE_2823));


OneBitAdder	b2v_inst963(
	.ci(SYNTHESIZED_WIRE_2829),
	.a(SYNTHESIZED_WIRE_2830),
	.b(SYNTHESIZED_WIRE_2831),
	.co(SYNTHESIZED_WIRE_2832),
	.s(SYNTHESIZED_WIRE_2724));


OneBitAdder	b2v_inst964(
	.ci(SYNTHESIZED_WIRE_2832),
	.a(SYNTHESIZED_WIRE_2833),
	.b(SYNTHESIZED_WIRE_2834),
	.co(SYNTHESIZED_WIRE_2835),
	.s(SYNTHESIZED_WIRE_2727));


OneBitAdder	b2v_inst965(
	.ci(SYNTHESIZED_WIRE_2835),
	.a(SYNTHESIZED_WIRE_2836),
	.b(SYNTHESIZED_WIRE_2837),
	.co(SYNTHESIZED_WIRE_2838),
	.s(SYNTHESIZED_WIRE_2730));


OneBitAdder	b2v_inst966(
	.ci(SYNTHESIZED_WIRE_2838),
	.a(SYNTHESIZED_WIRE_2839),
	.b(SYNTHESIZED_WIRE_2840),
	.co(SYNTHESIZED_WIRE_2841),
	.s(SYNTHESIZED_WIRE_2733));


OneBitAdder	b2v_inst967(
	.ci(SYNTHESIZED_WIRE_2841),
	.a(SYNTHESIZED_WIRE_2842),
	.b(SYNTHESIZED_WIRE_2843),
	.co(SYNTHESIZED_WIRE_2844),
	.s(SYNTHESIZED_WIRE_2736));


OneBitAdder	b2v_inst968(
	.ci(SYNTHESIZED_WIRE_2844),
	.a(SYNTHESIZED_WIRE_2845),
	.b(SYNTHESIZED_WIRE_2846),
	.co(SYNTHESIZED_WIRE_2847),
	.s(SYNTHESIZED_WIRE_2739));


OneBitAdder	b2v_inst969(
	.ci(SYNTHESIZED_WIRE_2847),
	.a(SYNTHESIZED_WIRE_2848),
	.b(SYNTHESIZED_WIRE_2849),
	.co(SYNTHESIZED_WIRE_2852),
	.s(SYNTHESIZED_WIRE_2742));


OneBitAdderHalf	b2v_inst97(
	.A(SYNTHESIZED_WIRE_2850),
	.B(SYNTHESIZED_WIRE_2851),
	.C(SYNTHESIZED_WIRE_116),
	.S(Z_ALTERA_SYNTHESIZED[29]));


OneBitAdder	b2v_inst970(
	.ci(SYNTHESIZED_WIRE_2852),
	.a(SYNTHESIZED_WIRE_2853),
	.b(SYNTHESIZED_WIRE_2854),
	.co(SYNTHESIZED_WIRE_2855),
	.s(SYNTHESIZED_WIRE_2745));


OneBitAdder	b2v_inst971(
	.ci(SYNTHESIZED_WIRE_2855),
	.a(SYNTHESIZED_WIRE_2856),
	.b(SYNTHESIZED_WIRE_2857),
	.co(SYNTHESIZED_WIRE_2858),
	.s(SYNTHESIZED_WIRE_2748));


OneBitAdder	b2v_inst972(
	.ci(SYNTHESIZED_WIRE_2858),
	.a(SYNTHESIZED_WIRE_2859),
	.b(SYNTHESIZED_WIRE_2860),
	.co(SYNTHESIZED_WIRE_2861),
	.s(SYNTHESIZED_WIRE_2751));


OneBitAdder	b2v_inst973(
	.ci(SYNTHESIZED_WIRE_2861),
	.a(SYNTHESIZED_WIRE_2862),
	.b(SYNTHESIZED_WIRE_2863),
	.co(SYNTHESIZED_WIRE_2864),
	.s(SYNTHESIZED_WIRE_2757));


OneBitAdder	b2v_inst974(
	.ci(SYNTHESIZED_WIRE_2864),
	.a(SYNTHESIZED_WIRE_2865),
	.b(SYNTHESIZED_WIRE_2866),
	.co(SYNTHESIZED_WIRE_2867),
	.s(SYNTHESIZED_WIRE_2760));


OneBitAdder	b2v_inst975(
	.ci(SYNTHESIZED_WIRE_2867),
	.a(SYNTHESIZED_WIRE_2868),
	.b(SYNTHESIZED_WIRE_2869),
	.co(SYNTHESIZED_WIRE_2870),
	.s(SYNTHESIZED_WIRE_2763));


OneBitAdder	b2v_inst976(
	.ci(SYNTHESIZED_WIRE_2870),
	.a(SYNTHESIZED_WIRE_2871),
	.b(SYNTHESIZED_WIRE_2872),
	.co(SYNTHESIZED_WIRE_2769),
	.s(SYNTHESIZED_WIRE_2766));


OneBitAdder	b2v_inst977(
	.ci(SYNTHESIZED_WIRE_2873),
	.a(SYNTHESIZED_WIRE_2874),
	.b(SYNTHESIZED_WIRE_2875),
	.co(SYNTHESIZED_WIRE_2876),
	.s(SYNTHESIZED_WIRE_2717));


OneBitAdder	b2v_inst978(
	.ci(SYNTHESIZED_WIRE_2876),
	.a(SYNTHESIZED_WIRE_2877),
	.b(SYNTHESIZED_WIRE_2878),
	.co(SYNTHESIZED_WIRE_2879),
	.s(SYNTHESIZED_WIRE_2772));


OneBitAdder	b2v_inst979(
	.ci(SYNTHESIZED_WIRE_2879),
	.a(SYNTHESIZED_WIRE_2880),
	.b(SYNTHESIZED_WIRE_2881),
	.co(SYNTHESIZED_WIRE_2885),
	.s(SYNTHESIZED_WIRE_2775));


OneBitAdder	b2v_inst98(
	.ci(SYNTHESIZED_WIRE_2882),
	.a(SYNTHESIZED_WIRE_2883),
	.b(SYNTHESIZED_WIRE_2884),
	.co(SYNTHESIZED_WIRE_2915),
	.s(SYNTHESIZED_WIRE_2820));


OneBitAdder	b2v_inst980(
	.ci(SYNTHESIZED_WIRE_2885),
	.a(SYNTHESIZED_WIRE_2886),
	.b(SYNTHESIZED_WIRE_2887),
	.co(SYNTHESIZED_WIRE_2888),
	.s(SYNTHESIZED_WIRE_2778));


OneBitAdder	b2v_inst981(
	.ci(SYNTHESIZED_WIRE_2888),
	.a(SYNTHESIZED_WIRE_2889),
	.b(SYNTHESIZED_WIRE_2890),
	.co(SYNTHESIZED_WIRE_2891),
	.s(SYNTHESIZED_WIRE_2781));


OneBitAdder	b2v_inst982(
	.ci(SYNTHESIZED_WIRE_2891),
	.a(SYNTHESIZED_WIRE_2892),
	.b(SYNTHESIZED_WIRE_2893),
	.co(SYNTHESIZED_WIRE_2894),
	.s(SYNTHESIZED_WIRE_2784));


OneBitAdder	b2v_inst983(
	.ci(SYNTHESIZED_WIRE_2894),
	.a(SYNTHESIZED_WIRE_2895),
	.b(SYNTHESIZED_WIRE_2896),
	.co(SYNTHESIZED_WIRE_2897),
	.s(SYNTHESIZED_WIRE_2790));


OneBitAdder	b2v_inst984(
	.ci(SYNTHESIZED_WIRE_2897),
	.a(SYNTHESIZED_WIRE_2898),
	.b(SYNTHESIZED_WIRE_2899),
	.co(SYNTHESIZED_WIRE_2900),
	.s(SYNTHESIZED_WIRE_2793));


OneBitAdder	b2v_inst985(
	.ci(SYNTHESIZED_WIRE_2900),
	.a(SYNTHESIZED_WIRE_2901),
	.b(SYNTHESIZED_WIRE_2902),
	.co(SYNTHESIZED_WIRE_2903),
	.s(SYNTHESIZED_WIRE_2796));


OneBitAdder	b2v_inst986(
	.ci(SYNTHESIZED_WIRE_2903),
	.a(SYNTHESIZED_WIRE_2904),
	.b(SYNTHESIZED_WIRE_2905),
	.co(SYNTHESIZED_WIRE_2906),
	.s(SYNTHESIZED_WIRE_2799));


OneBitAdder	b2v_inst987(
	.ci(SYNTHESIZED_WIRE_2906),
	.a(SYNTHESIZED_WIRE_2907),
	.b(SYNTHESIZED_WIRE_2908),
	.co(SYNTHESIZED_WIRE_2909),
	.s(SYNTHESIZED_WIRE_2802));


OneBitAdder	b2v_inst988(
	.ci(SYNTHESIZED_WIRE_2909),
	.a(SYNTHESIZED_WIRE_2910),
	.b(SYNTHESIZED_WIRE_2911),
	.co(SYNTHESIZED_WIRE_2912),
	.s(SYNTHESIZED_WIRE_2805));


OneBitAdder	b2v_inst989(
	.ci(SYNTHESIZED_WIRE_2912),
	.a(SYNTHESIZED_WIRE_2913),
	.b(SYNTHESIZED_WIRE_2914),
	.co(SYNTHESIZED_WIRE_2918),
	.s(SYNTHESIZED_WIRE_2808));


OneBitAdder	b2v_inst99(
	.ci(SYNTHESIZED_WIRE_2915),
	.a(SYNTHESIZED_WIRE_2916),
	.b(SYNTHESIZED_WIRE_2917),
	.co(SYNTHESIZED_WIRE_2),
	.s(SYNTHESIZED_WIRE_1839));


OneBitAdder	b2v_inst990(
	.ci(SYNTHESIZED_WIRE_2918),
	.a(SYNTHESIZED_WIRE_2919),
	.b(SYNTHESIZED_WIRE_2920),
	.co(SYNTHESIZED_WIRE_2921),
	.s(SYNTHESIZED_WIRE_2811));


OneBitAdder	b2v_inst991(
	.ci(SYNTHESIZED_WIRE_2921),
	.a(SYNTHESIZED_WIRE_2922),
	.b(SYNTHESIZED_WIRE_2923),
	.co(SYNTHESIZED_WIRE_2924),
	.s(SYNTHESIZED_WIRE_2814));


OneBitAdder	b2v_inst992(
	.ci(SYNTHESIZED_WIRE_2924),
	.a(SYNTHESIZED_WIRE_2925),
	.b(SYNTHESIZED_WIRE_2926),
	.co(SYNTHESIZED_WIRE_2826),
	.s(SYNTHESIZED_WIRE_2817));


OneBitAdderHalf	b2v_inst993(
	.A(SYNTHESIZED_WIRE_2927),
	.B(SYNTHESIZED_WIRE_2928),
	.C(SYNTHESIZED_WIRE_32),
	.S(Z_ALTERA_SYNTHESIZED[1]));


OneBitAdder	b2v_inst994(
	.ci(SYNTHESIZED_WIRE_2929),
	.a(SYNTHESIZED_WIRE_2930),
	.b(SYNTHESIZED_WIRE_2931),
	.co(SYNTHESIZED_WIRE_2932),
	.s(SYNTHESIZED_WIRE_2926));


OneBitAdder	b2v_inst995(
	.ci(SYNTHESIZED_WIRE_2932),
	.a(SYNTHESIZED_WIRE_2933),
	.b(SYNTHESIZED_WIRE_2934),
	.co(SYNTHESIZED_WIRE_2935),
	.s(SYNTHESIZED_WIRE_2828));


OneBitAdder	b2v_inst996(
	.ci(SYNTHESIZED_WIRE_2935),
	.a(SYNTHESIZED_WIRE_2936),
	.b(SYNTHESIZED_WIRE_2937),
	.co(SYNTHESIZED_WIRE_2938),
	.s(SYNTHESIZED_WIRE_2831));


OneBitAdder	b2v_inst997(
	.ci(SYNTHESIZED_WIRE_2938),
	.a(SYNTHESIZED_WIRE_2939),
	.b(SYNTHESIZED_WIRE_2940),
	.co(SYNTHESIZED_WIRE_2941),
	.s(SYNTHESIZED_WIRE_2834));


OneBitAdder	b2v_inst998(
	.ci(SYNTHESIZED_WIRE_2941),
	.a(SYNTHESIZED_WIRE_2942),
	.b(SYNTHESIZED_WIRE_2943),
	.co(SYNTHESIZED_WIRE_2944),
	.s(SYNTHESIZED_WIRE_2837));


OneBitAdder	b2v_inst999(
	.ci(SYNTHESIZED_WIRE_2944),
	.a(SYNTHESIZED_WIRE_2945),
	.b(SYNTHESIZED_WIRE_2946),
	.co(SYNTHESIZED_WIRE_5),
	.s(SYNTHESIZED_WIRE_2840));

assign	Z = Z_ALTERA_SYNTHESIZED;

endmodule
