///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: SE16_32
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();
`include "../Test/Test.v"
///////////////////////////////////////////////////////////////////////////////////
// Input: A, B (32-bit) 
reg[31:0] A, B;
///////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
// Output: Z (64-bit)
wire[63:0] Z;
///////////////////////////////////////////////////////////////////////////////////

Multiplier_32 myMultiplier(.A(A), .B(B), .Z(Z));

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: Two positives
$display("Testing two positives: 14*3=42");
A=14;  B=3;   #10; 
verifyEqual64(Z, 42);
////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////
// Test: Positive-negative
$display("Testing positive-negative: 100*-20=2000");
A=100; B=-20;  #10;
verifyEqual64(Z, -2000);
////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////
// Test: Negative-positive
$display("Testing negative-positive: -75*4=-300");
A=-75;  B=4;   #10; 
verifyEqual64(Z, -300);
////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////
// Test: Two negatives
$display("Testing two negatives: -55*-10=550");
A=-55; B=-10;  #10;
verifyEqual64(Z, 550);
////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////
// Test: Multiplication by zero
$display("Testing multiplication by zero: 289*0=0");
A=289; B=0;  #10;
verifyEqual64(Z, 0);
////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////
// Test: Multiplication by one
$display("Testing multiplication by one: 1*-3817=-3817");
A=1; B=-3817;  #10;
verifyEqual64(Z, -3817);
////////////////////////////////////////////////////////////////////////////////////////

$display("All tests passed.");
end

endmodule